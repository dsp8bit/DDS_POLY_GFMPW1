VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DDS_Module
  CLASS BLOCK ;
  FOREIGN DDS_Module ;
  ORIGIN 0.000 0.000 ;
  SIZE 629.660 BY 647.580 ;
  PIN Cos_Out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 228.480 629.660 229.040 ;
    END
  END Cos_Out[0]
  PIN Cos_Out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 497.280 629.660 497.840 ;
    END
  END Cos_Out[10]
  PIN Cos_Out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 524.160 629.660 524.720 ;
    END
  END Cos_Out[11]
  PIN Cos_Out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 551.040 629.660 551.600 ;
    END
  END Cos_Out[12]
  PIN Cos_Out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 577.920 629.660 578.480 ;
    END
  END Cos_Out[13]
  PIN Cos_Out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 604.800 629.660 605.360 ;
    END
  END Cos_Out[14]
  PIN Cos_Out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 631.680 629.660 632.240 ;
    END
  END Cos_Out[15]
  PIN Cos_Out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 255.360 629.660 255.920 ;
    END
  END Cos_Out[1]
  PIN Cos_Out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 282.240 629.660 282.800 ;
    END
  END Cos_Out[2]
  PIN Cos_Out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 309.120 629.660 309.680 ;
    END
  END Cos_Out[3]
  PIN Cos_Out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 336.000 629.660 336.560 ;
    END
  END Cos_Out[4]
  PIN Cos_Out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 362.880 629.660 363.440 ;
    END
  END Cos_Out[5]
  PIN Cos_Out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 389.760 629.660 390.320 ;
    END
  END Cos_Out[6]
  PIN Cos_Out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 416.640 629.660 417.200 ;
    END
  END Cos_Out[7]
  PIN Cos_Out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 443.520 629.660 444.080 ;
    END
  END Cos_Out[8]
  PIN Cos_Out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 470.400 629.660 470.960 ;
    END
  END Cos_Out[9]
  PIN Enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END Enable
  PIN FreqPhase[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END FreqPhase[0]
  PIN FreqPhase[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END FreqPhase[10]
  PIN FreqPhase[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 488.320 0.000 488.880 4.000 ;
    END
  END FreqPhase[11]
  PIN FreqPhase[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 0.000 518.000 4.000 ;
    END
  END FreqPhase[12]
  PIN FreqPhase[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 546.560 0.000 547.120 4.000 ;
    END
  END FreqPhase[13]
  PIN FreqPhase[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 0.000 576.240 4.000 ;
    END
  END FreqPhase[14]
  PIN FreqPhase[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 0.000 605.360 4.000 ;
    END
  END FreqPhase[15]
  PIN FreqPhase[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 0.000 197.680 4.000 ;
    END
  END FreqPhase[1]
  PIN FreqPhase[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END FreqPhase[2]
  PIN FreqPhase[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END FreqPhase[3]
  PIN FreqPhase[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END FreqPhase[4]
  PIN FreqPhase[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 0.000 314.160 4.000 ;
    END
  END FreqPhase[5]
  PIN FreqPhase[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 0.000 343.280 4.000 ;
    END
  END FreqPhase[6]
  PIN FreqPhase[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 371.840 0.000 372.400 4.000 ;
    END
  END FreqPhase[7]
  PIN FreqPhase[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 0.000 401.520 4.000 ;
    END
  END FreqPhase[8]
  PIN FreqPhase[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 0.000 430.640 4.000 ;
    END
  END FreqPhase[9]
  PIN LoadF
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END LoadF
  PIN LoadP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 0.000 110.320 4.000 ;
    END
  END LoadP
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 0.000 22.960 4.000 ;
    END
  END clk
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 13.440 629.660 14.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 443.520 4.000 444.080 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.880 4.000 363.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 282.240 4.000 282.800 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 4.000 40.880 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 40.320 629.660 40.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 67.200 629.660 67.760 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 94.080 629.660 94.640 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 120.960 629.660 121.520 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 147.840 629.660 148.400 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 174.720 629.660 175.280 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 625.660 201.600 629.660 202.160 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 604.800 4.000 605.360 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 524.160 4.000 524.720 ;
    END
  END io_oeb[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 631.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 631.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 631.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 631.420 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 631.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 631.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 631.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 631.420 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 622.720 631.420 ;
      LAYER Metal2 ;
        RECT 6.300 4.300 622.020 632.150 ;
        RECT 6.300 3.500 22.100 4.300 ;
        RECT 23.260 3.500 51.220 4.300 ;
        RECT 52.380 3.500 80.340 4.300 ;
        RECT 81.500 3.500 109.460 4.300 ;
        RECT 110.620 3.500 138.580 4.300 ;
        RECT 139.740 3.500 167.700 4.300 ;
        RECT 168.860 3.500 196.820 4.300 ;
        RECT 197.980 3.500 225.940 4.300 ;
        RECT 227.100 3.500 255.060 4.300 ;
        RECT 256.220 3.500 284.180 4.300 ;
        RECT 285.340 3.500 313.300 4.300 ;
        RECT 314.460 3.500 342.420 4.300 ;
        RECT 343.580 3.500 371.540 4.300 ;
        RECT 372.700 3.500 400.660 4.300 ;
        RECT 401.820 3.500 429.780 4.300 ;
        RECT 430.940 3.500 458.900 4.300 ;
        RECT 460.060 3.500 488.020 4.300 ;
        RECT 489.180 3.500 517.140 4.300 ;
        RECT 518.300 3.500 546.260 4.300 ;
        RECT 547.420 3.500 575.380 4.300 ;
        RECT 576.540 3.500 604.500 4.300 ;
        RECT 605.660 3.500 622.020 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 631.380 625.360 632.100 ;
        RECT 4.000 605.660 625.660 631.380 ;
        RECT 4.300 604.500 625.360 605.660 ;
        RECT 4.000 578.780 625.660 604.500 ;
        RECT 4.000 577.620 625.360 578.780 ;
        RECT 4.000 551.900 625.660 577.620 ;
        RECT 4.000 550.740 625.360 551.900 ;
        RECT 4.000 525.020 625.660 550.740 ;
        RECT 4.300 523.860 625.360 525.020 ;
        RECT 4.000 498.140 625.660 523.860 ;
        RECT 4.000 496.980 625.360 498.140 ;
        RECT 4.000 471.260 625.660 496.980 ;
        RECT 4.000 470.100 625.360 471.260 ;
        RECT 4.000 444.380 625.660 470.100 ;
        RECT 4.300 443.220 625.360 444.380 ;
        RECT 4.000 417.500 625.660 443.220 ;
        RECT 4.000 416.340 625.360 417.500 ;
        RECT 4.000 390.620 625.660 416.340 ;
        RECT 4.000 389.460 625.360 390.620 ;
        RECT 4.000 363.740 625.660 389.460 ;
        RECT 4.300 362.580 625.360 363.740 ;
        RECT 4.000 336.860 625.660 362.580 ;
        RECT 4.000 335.700 625.360 336.860 ;
        RECT 4.000 309.980 625.660 335.700 ;
        RECT 4.000 308.820 625.360 309.980 ;
        RECT 4.000 283.100 625.660 308.820 ;
        RECT 4.300 281.940 625.360 283.100 ;
        RECT 4.000 256.220 625.660 281.940 ;
        RECT 4.000 255.060 625.360 256.220 ;
        RECT 4.000 229.340 625.660 255.060 ;
        RECT 4.000 228.180 625.360 229.340 ;
        RECT 4.000 202.460 625.660 228.180 ;
        RECT 4.300 201.300 625.360 202.460 ;
        RECT 4.000 175.580 625.660 201.300 ;
        RECT 4.000 174.420 625.360 175.580 ;
        RECT 4.000 148.700 625.660 174.420 ;
        RECT 4.000 147.540 625.360 148.700 ;
        RECT 4.000 121.820 625.660 147.540 ;
        RECT 4.300 120.660 625.360 121.820 ;
        RECT 4.000 94.940 625.660 120.660 ;
        RECT 4.000 93.780 625.360 94.940 ;
        RECT 4.000 68.060 625.660 93.780 ;
        RECT 4.000 66.900 625.360 68.060 ;
        RECT 4.000 41.180 625.660 66.900 ;
        RECT 4.300 40.020 625.360 41.180 ;
        RECT 4.000 14.300 625.660 40.020 ;
        RECT 4.000 13.580 625.360 14.300 ;
      LAYER Metal4 ;
        RECT 16.380 27.530 21.940 596.870 ;
        RECT 24.140 27.530 98.740 596.870 ;
        RECT 100.940 27.530 175.540 596.870 ;
        RECT 177.740 27.530 252.340 596.870 ;
        RECT 254.540 27.530 329.140 596.870 ;
        RECT 331.340 27.530 405.940 596.870 ;
        RECT 408.140 27.530 482.740 596.870 ;
        RECT 484.940 27.530 559.540 596.870 ;
        RECT 561.740 27.530 602.420 596.870 ;
  END
END DDS_Module
END LIBRARY

