// This is the unpowered netlist.
module DDS_Module (Enable,
    LoadF,
    LoadP,
    clk,
    rst,
    Cos_Out,
    FreqPhase,
    io_oeb);
 input Enable;
 input LoadF;
 input LoadP;
 input clk;
 input rst;
 output [15:0] Cos_Out;
 input [15:0] FreqPhase;
 output [15:0] io_oeb;

 wire net37;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-10] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-11] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-12] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-13] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-14] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-15] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-16] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-17] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-18] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-19] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-20] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-21] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-22] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-23] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-24] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-25] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-5] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-6] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-7] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-8] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-9] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[0] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-10] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-11] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-12] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-13] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-14] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-15] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-16] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-17] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-18] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-19] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-20] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-21] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-22] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-23] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-24] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-25] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-6] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-7] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-8] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[5] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-10] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-11] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-12] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-13] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-14] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-15] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-16] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-17] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-18] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-19] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-20] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-21] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-22] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-23] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-24] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-25] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-5] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-6] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-7] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-8] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-9] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[0] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[5] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-10] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-11] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-12] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-13] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-14] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-15] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-16] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-17] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-18] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-19] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-20] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-21] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-22] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-23] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-24] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-25] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-5] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-6] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-7] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-8] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-9] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[0] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-10] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-11] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-12] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-13] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-14] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-15] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-5] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-6] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-7] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-8] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-9] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-10] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-11] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-12] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-13] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-14] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-15] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-5] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-6] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-7] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-8] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-9] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[0] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[10] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[11] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[12] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[13] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[14] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[15] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[16] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[17] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[18] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[19] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[20] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[21] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[22] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[23] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[24] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[25] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[26] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[27] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[28] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[29] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[30] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[31] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[5] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[6] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[7] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[8] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[9] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[0] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[1] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[2] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[3] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[4] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[16] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[17] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[18] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[19] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[20] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[21] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[22] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[23] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[24] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[25] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[26] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[27] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[28] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[29] ;
 wire \DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[30] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-10] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-11] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-12] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-14] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-15] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-1] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-2] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-3] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-4] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-5] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-6] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-7] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-8] ;
 wire \DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-9] ;
 wire \DDS_Stage.LCU.SelMuxConfig ;
 wire \DDS_Stage.LCU.SelMuxConfigReg ;
 wire \DDS_Stage.LCU.state[0] ;
 wire \DDS_Stage.LCU.state[1] ;
 wire \DDS_Stage.LCU.state[2] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-10] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-11] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-12] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-13] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-14] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-15] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-1] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-2] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-3] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-4] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-5] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-6] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-7] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-8] ;
 wire \DDS_Stage.xPoints_Generator1.CosNew[-9] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-10] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-11] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-12] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-13] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-14] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-15] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-1] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-2] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-3] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-4] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-5] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-6] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-7] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-8] ;
 wire \DDS_Stage.xPoints_Generator1.RegF[-9] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-10] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-11] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-12] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-13] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-14] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-15] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-1] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-2] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-3] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-4] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-5] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-6] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-7] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-8] ;
 wire \DDS_Stage.xPoints_Generator1.RegFrequency[-9] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-10] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-11] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-12] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-13] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-14] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-15] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-1] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-2] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-3] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-4] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-5] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-6] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-7] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-8] ;
 wire \DDS_Stage.xPoints_Generator1.RegP[-9] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net4;
 wire net5;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__I (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__I (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__I (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__I (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__I (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A1 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__A1 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__A2 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__A1 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__A2 (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A2 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__I (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A2 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A2 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__A2 (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A1 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__I (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A1 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A2 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__A2 (.I(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A2 (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A2 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A2 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__I (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A1 (.I(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A2 (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A1 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__A2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__A1 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__A2 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A1 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__A2 (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__B (.I(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__C (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__B (.I(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06915__I0 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06915__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__I (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__A1 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__B (.I(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__A2 (.I(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__B2 (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__A2 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A2 (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__I (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A2 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A2 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__I (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A2 (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A2 (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06942__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06946__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06946__A2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06946__B (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A1 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A2 (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A2 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A3 (.I(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__A2 (.I(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A2 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A2 (.I(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__B2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__A2 (.I(_06576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__A2 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A2 (.I(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__B (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__C (.I(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A2 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__A1 (.I(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A2 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A2 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A2 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A1 (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A2 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A2 (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A3 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__B (.I(_06646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__A2 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A2 (.I(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A3 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__A2 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A1 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A2 (.I(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A1 (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A2 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A2 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__A1 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A2 (.I(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__A2 (.I(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__A1 (.I(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07056__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__A2 (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__A2 (.I(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A2 (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__B2 (.I(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__A2 (.I(_06700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07077__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07077__A2 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__B (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A2 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__A1 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__I0 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A2 (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__B (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A1 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A2 (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__A2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__B (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A1 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A1 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A2 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07112__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07112__A2 (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A2 (.I(_06732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__A2 (.I(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A1 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A2 (.I(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__B (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07119__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A2 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A2 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__B (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A1 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A1 (.I(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__A2 (.I(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__A2 (.I(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__A2 (.I(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__B (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__A2 (.I(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07144__B (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__A2 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__B (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__A2 (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A2 (.I(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__A2 (.I(_06732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07156__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__A1 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__A2 (.I(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07163__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07163__A2 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__C (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A2 (.I(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__B (.I(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A1 (.I(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A2 (.I(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__B (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A2 (.I(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__B (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A1 (.I(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A2 (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__B (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__A1 (.I(_06787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A2 (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A3 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A4 (.I(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A1 (.I(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__A2 (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__B (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A2 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__B1 (.I(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__I1 (.I(_06800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__A2 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A2 (.I(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__I1 (.I(_06804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__A2 (.I(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__B2 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A2 (.I(_06809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__A1 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__B1 (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__B2 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__A2 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A1 (.I(_06646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A2 (.I(_06811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__B2 (.I(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__I1 (.I(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A3 (.I(_06787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A1 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A2 (.I(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__B2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__B2 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__C (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__B (.I(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__A2 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__B1 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__B2 (.I(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__B (.I(_06829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A3 (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A2 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A3 (.I(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A2 (.I(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A2 (.I(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A2 (.I(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A2 (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A2 (.I(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A1 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__B (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__C (.I(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A2 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A3 (.I(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A1 (.I(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A2 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A1 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__B (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__A2 (.I(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A2 (.I(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__C (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A1 (.I(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A1 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A2 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__B1 (.I(_06732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__B2 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A2 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__I1 (.I(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__B1 (.I(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__B2 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__A2 (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A2 (.I(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__B1 (.I(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A2 (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__B2 (.I(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__C (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A3 (.I(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__A2 (.I(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A2 (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A2 (.I(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__C (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__B (.I(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A1 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__B1 (.I(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__B2 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A2 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A1 (.I(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A2 (.I(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A2 (.I(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A2 (.I(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A1 (.I(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__B (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__B (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A1 (.I(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A2 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__B (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__I0 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__I1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__I0 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__I1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A2 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__A2 (.I(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__I0 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__I1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__I0 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__I1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__I0 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__I1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__I0 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__I1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__I0 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__I1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__I0 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__I1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__I0 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__I1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__I0 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__I1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__I0 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__I1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__I0 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__I1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__S (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__I (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__I0 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__I1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__I0 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__I1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A2 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__C (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A1 (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A2 (.I(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__A1 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A1 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__C (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__B (.I(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A2 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__B (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__A2 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__B (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A2 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__B2 (.I(_06732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A2 (.I(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A1 (.I(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__B2 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A2 (.I(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A1 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A2 (.I(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A1 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__C (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__B (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__C (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A2 (.I(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__B (.I(_06646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A2 (.I(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A1 (.I(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__B2 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A2 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A3 (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__B (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__B1 (.I(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A2 (.I(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A1 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A2 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__B2 (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A2 (.I(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A1 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__B2 (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__A1 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A2 (.I(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__C (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A1 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A2 (.I(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__B (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A2 (.I(_06787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A2 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A3 (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__B (.I(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A1 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__B2 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__C (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A1 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A2 (.I(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A2 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A1 (.I(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__B2 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A1 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A2 (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__B1 (.I(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__B2 (.I(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__A2 (.I(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__B2 (.I(_06787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A1 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__B (.I(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__A2 (.I(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A2 (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A3 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A1 (.I(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A1 (.I(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__B (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__B (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A2 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__B1 (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A2 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A3 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A2 (.I(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A3 (.I(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__A1 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A2 (.I(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__B (.I(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A1 (.I(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__B (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__C (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A2 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A2 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A1 (.I(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A2 (.I(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A2 (.I(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A2 (.I(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__B1 (.I(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A2 (.I(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A2 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__C (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__B (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A1 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__A1 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__B (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A2 (.I(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A3 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A2 (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__B (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A1 (.I(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__B2 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__I0 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A1 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A2 (.I(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__B (.I(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A2 (.I(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A2 (.I(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__B1 (.I(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A2 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__C (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A1 (.I(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A1 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A2 (.I(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__A3 (.I(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__A1 (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A2 (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__A2 (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__A1 (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__I0 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__I1 (.I(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A2 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__B (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__A2 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__B (.I(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A2 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__B (.I(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__A2 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__B (.I(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A2 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__B (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__I (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A2 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__A2 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A1 (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__A1 (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A1 (.I(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__I0 (.I(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A1 (.I(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A1 (.I(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__S (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__I0 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__S (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__S (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__S (.I(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__I0 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__I0 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A2 (.I(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__B (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__I0 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__I0 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__I (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__I0 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__I0 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__I0 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__I0 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__I0 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A2 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A1 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A1 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A3 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A4 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A1 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__B1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__B2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A3 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A4 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A1 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__B1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__B2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A1 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A3 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A4 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A1 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A3 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A4 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A2 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__B1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__B2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A2 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__B1 (.I(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__B2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A3 (.I(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A4 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A1 (.I(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A2 (.I(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__B1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__B2 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A3 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A4 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A2 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__B1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__B2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A3 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A4 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__B1 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__B2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A3 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A4 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A2 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A1 (.I(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A2 (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A1 (.I(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A1 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A3 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A4 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A3 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A4 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__B1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__B2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__B1 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__B2 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A3 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A4 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A2 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A2 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A2 (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A3 (.I(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A4 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__A2 (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__B1 (.I(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__B2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A2 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__B1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__B2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A2 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A3 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A4 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A2 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A2 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A2 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A2 (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A3 (.I(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A4 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A2 (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__B1 (.I(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__B2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A1 (.I(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A1 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A1 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A1 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__B1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__B2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A1 (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A2 (.I(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__B1 (.I(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__B2 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A3 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A4 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A2 (.I(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A1 (.I(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A2 (.I(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A1 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A3 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A4 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A1 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__B1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__B2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A3 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A4 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__B1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__B2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__B1 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__B2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A3 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A4 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A2 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__B1 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__B2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A3 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A4 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__B1 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__B2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A3 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A4 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A2 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__B1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__B2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A3 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A4 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A2 (.I(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A1 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A3 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__A4 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__B1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__B2 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A3 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A4 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A2 (.I(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A1 (.I(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A1 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A3 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A4 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A1 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__B1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__B2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A1 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A2 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A3 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A4 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A3 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A4 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__B1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__B2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__B1 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A1 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A3 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A4 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__B (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__C (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A1 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A1 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A2 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A2 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A1 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A1 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A2 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__B1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__B2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A3 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A4 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A2 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A1 (.I(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A2 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A2 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A1 (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A2 (.I(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A1 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A2 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A2 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__I0 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A2 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__A1 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A2 (.I(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A2 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A2 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__B2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A3 (.I(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A4 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A3 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A4 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__B1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__B2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__B1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__B2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A3 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A4 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A2 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A2 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__B2 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__A2 (.I(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A3 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A4 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A1 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__B2 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A2 (.I(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A3 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A4 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__B1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__B2 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A3 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A4 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A2 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A2 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A3 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A4 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A2 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__B1 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__B2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A2 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A2 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A3 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A4 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__B2 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A1 (.I(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A3 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A4 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A2 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A2 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__B1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A3 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A4 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A2 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A2 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__B1 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__B2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A3 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A4 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A2 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A2 (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A2 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__B1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A3 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A4 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A1 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A2 (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A1 (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A2 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__B1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__B2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A3 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A4 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A2 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A2 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__B1 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A3 (.I(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__A4 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__B1 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__B2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A3 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A4 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A2 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A2 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__B1 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__B2 (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A3 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A4 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__B1 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__B2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A3 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A4 (.I(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A1 (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A2 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__B1 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A3 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A4 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A2 (.I(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A2 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A2 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__B1 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__B2 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A3 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A4 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__B1 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A3 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A4 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__A2 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A2 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A2 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A2 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A2 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A1 (.I(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__B1 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A3 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A4 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A1 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A2 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__A2 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A2 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__A1 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__B2 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A2 (.I(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A3 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A4 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__B1 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A3 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A4 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09344__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__B1 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__B2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A3 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A4 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__B1 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__B2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A3 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A4 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__B2 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A2 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A3 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A4 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__I0 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__I1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__B1 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__B2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A3 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A4 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__B1 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__B2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A3 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A4 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A1 (.I(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A2 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A2 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A1 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A2 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__B1 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__B2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A3 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A4 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__B2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A1 (.I(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A3 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A4 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A1 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A2 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__B1 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__B2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A3 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A4 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A1 (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__B2 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A3 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A4 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__B1 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__B2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A2 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A3 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A4 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A1 (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A1 (.I(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A1 (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A1 (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__B1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__B2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A1 (.I(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A2 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A3 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A4 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__I0 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__I1 (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A1 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A1 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__B1 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A3 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A4 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A1 (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A3 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__B (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A3 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__B1 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A3 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A4 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__I (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__B1 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A3 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A4 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__B (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A3 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A2 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__B1 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A3 (.I(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A4 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A3 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A4 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__B1 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__B2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A1 (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A1 (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__B1 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__B2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A3 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A4 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__B (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A3 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__A2 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__B1 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A3 (.I(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A4 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__B (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A3 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A2 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__B1 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A3 (.I(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A4 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__I0 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__I1 (.I(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__S (.I(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A1 (.I(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__B (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__B (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__B (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__B (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A3 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A2 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__B1 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A3 (.I(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A4 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A1 (.I(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A2 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__B (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A2 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A4 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__B (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A3 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A2 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__B1 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A3 (.I(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A4 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A1 (.I(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A1 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__B (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A3 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A2 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__B1 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A3 (.I(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A4 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A1 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A2 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A2 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__B (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A3 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A2 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__B1 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A3 (.I(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A4 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__B (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A2 (.I(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A3 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A2 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A2 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__B (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__A3 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__A2 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__B1 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A3 (.I(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A4 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A2 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__A2 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__B (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A3 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A2 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__B1 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A3 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A4 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__A1 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__A1 (.I(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__B (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A3 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A2 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__B1 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__A3 (.I(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__A4 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__B (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A1 (.I(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A2 (.I(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A3 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__B2 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__B2 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A2 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__B (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A3 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A2 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__B1 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__B2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A3 (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A4 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A1 (.I(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__I0 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A1 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A2 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__B (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A2 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A3 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A1 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A1 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__B (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A1 (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__A2 (.I(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__B (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A1 (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A2 (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A2 (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__A1 (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__A1 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__A1 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A1 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A2 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__I0 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__I0 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__I0 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__I1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A2 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A2 (.I(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A2 (.I(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__I0 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__B (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A2 (.I(_06811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__I1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__I0 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A2 (.I(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__I0 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A3 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A4 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__B1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A3 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A4 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__B1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A3 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A4 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__B1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__B1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A3 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A4 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A2 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A2 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__B1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A3 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A4 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__A2 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A2 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A3 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A4 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__B1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A2 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__B1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A3 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A4 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A2 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A2 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A3 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A4 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__B1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__A2 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__B1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A3 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A4 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A2 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__B1 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__B2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A3 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A4 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__A2 (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A2 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A2 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__A2 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A2 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__B1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A3 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A4 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A3 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A4 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__B1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__B1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__B2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A3 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A4 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A2 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__B1 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A3 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A4 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A3 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A4 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A3 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A4 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__B1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__B1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A3 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A4 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A3 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A4 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__B1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A3 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A4 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__B1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__B2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__B1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A3 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A4 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__B1 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A3 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A4 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A1 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A1 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__B1 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A3 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A4 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__B1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A3 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A4 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__B1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__B2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A3 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A4 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11489__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11489__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__B1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A3 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A4 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__B1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A3 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A4 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A3 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A4 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__B1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11583__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11583__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11585__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11585__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__B1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A3 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A4 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__A3 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__A4 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11625__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11625__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__B1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A3 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A4 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11631__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11631__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__B1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__B2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__B1 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A3 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A4 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11647__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11647__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__A1 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__A3 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__A4 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__B1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__B2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11684__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11684__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11689__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11689__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11696__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11696__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__B1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__A3 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__A4 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11702__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11702__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11704__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11704__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__B1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__A3 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__A4 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__A3 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__A4 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__B1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__B2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11732__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11732__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__A3 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__A4 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__B1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__B2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11775__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11775__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__B1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__A3 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__A4 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11786__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11786__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11787__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11787__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__A3 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__A4 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11804__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11804__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__B1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__B2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11809__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11809__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__B1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__A3 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__A4 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11819__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11819__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__A3 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__A4 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__B1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__B2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11838__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11838__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11838__B1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11838__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__A3 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__A4 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11841__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11841__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11843__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11843__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11862__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11862__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__B1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11866__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11866__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11867__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11867__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11867__A3 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11867__A4 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11871__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11871__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11877__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11877__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__A3 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__A4 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11880__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11880__A2 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11895__A1 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11896__A1 (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11897__B1 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11899__A1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11899__A2 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11900__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11900__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__B1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11902__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11902__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11902__A3 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11902__A4 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11906__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11906__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11906__A3 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11906__A4 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__B1 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11911__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11911__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11913__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11913__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__A3 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__A4 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11918__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11918__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__B1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11923__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11923__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11925__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11925__A2 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__A3 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__A4 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__B1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11937__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11937__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11937__A3 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11937__A4 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__A3 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__A4 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11944__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11944__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11945__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11945__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11946__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11946__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__B1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__A3 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__A4 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11966__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11966__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11967__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11967__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11968__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11968__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11974__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11974__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11975__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11975__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11977__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11977__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11977__B1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11977__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__A3 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__A4 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11980__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11980__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11981__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11981__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12001__A2 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__A2 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12030__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12030__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__B1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__A3 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__A4 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__A3 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__A4 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12041__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12041__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__A3 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__A4 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12046__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12046__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__B1 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12051__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12051__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12052__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12052__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12053__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12053__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12074__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12074__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12075__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12075__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12075__B1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12075__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__A2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__A3 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__A4 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12078__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12078__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12100__A1 (.I(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12100__A2 (.I(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12102__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12102__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12103__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12103__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12103__B1 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12103__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__A3 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__A4 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__A3 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__A4 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12111__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12111__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12112__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12112__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12113__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12113__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12117__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12117__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12117__A3 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12117__A4 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12118__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12118__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12119__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12119__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12119__B1 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12119__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12124__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12124__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12125__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12125__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12147__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12147__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12148__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12148__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12148__B1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12148__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12149__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12149__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12149__A3 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12149__A4 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12151__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12151__A2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12152__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12152__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12178__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12178__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12179__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12179__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12179__A3 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12179__A4 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__B1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__B2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12184__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12184__A2 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12186__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12186__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12198__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12198__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12199__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12199__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12199__A3 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12199__A4 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__B1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__B2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__A3 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__A4 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__A3 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__A4 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12213__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12213__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12214__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12214__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__B1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__B2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__A2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__A3 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__A4 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12232__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12232__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__A1 (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12236__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12236__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12237__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12237__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12238__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12238__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12326__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12326__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12384__A1 (.I(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12384__A2 (.I(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12387__A1 (.I(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12387__A2 (.I(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12422__A1 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12437__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12437__B2 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12439__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12439__A2 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12441__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12442__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12442__A2 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__A2 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__B (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12446__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12446__A2 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12448__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12449__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12454__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12455__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12456__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12457__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__B2 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12477__A1 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12481__A1 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__A1 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12492__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12500__A1 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12506__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12506__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12516__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12516__A2 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12516__B1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12516__B2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12517__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12517__A2 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12517__A3 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12517__A4 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12519__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12519__A2 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__A2 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12521__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12521__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12524__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12524__A2 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__A1 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__A2 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12536__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12536__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12537__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12537__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12538__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12538__A2 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12548__A1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12548__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12549__A1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12549__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12550__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12550__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12556__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12556__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12557__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12557__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12558__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12558__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12578__A1 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12582__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12583__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12592__A1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12592__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__B1 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__B2 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__A2 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__A3 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__A4 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12605__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12605__A2 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12606__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12606__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12607__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12607__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12610__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12610__A2 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12611__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12611__A2 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12611__A3 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12611__A4 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__A2 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__B1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__B2 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12624__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12624__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12625__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12625__A2 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__A1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12638__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12638__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12639__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12639__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12645__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12645__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12646__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12646__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12647__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12647__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12667__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12668__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12669__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12677__A1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12677__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__A1 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__B1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__B2 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12687__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12687__A2 (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12687__A3 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12687__A4 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12689__A1 (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12689__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12690__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12690__A2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12690__A3 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12690__A4 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12691__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12691__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12691__B1 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12691__B2 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12694__A1 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12694__A2 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12695__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12695__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12696__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12696__A2 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12701__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12701__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12706__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12706__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__A2 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12719__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12719__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12720__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12720__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12721__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12721__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12727__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12727__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12728__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12728__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12729__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12729__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12758__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12767__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12767__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12781__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12781__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12782__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12782__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12783__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12783__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12786__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12786__A2 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12787__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12787__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12788__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12788__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12793__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12793__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12797__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12797__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12798__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12798__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12799__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12799__A2 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12814__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12814__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12815__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12815__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12822__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12822__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12823__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12823__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12824__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12824__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12842__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12843__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12844__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12859__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12859__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__B1 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__B2 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12870__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12870__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12870__A3 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12870__A4 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12873__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12873__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12873__B (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12874__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12874__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12874__A3 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12876__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12876__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12879__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12879__A2 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12880__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12880__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12892__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12892__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12893__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12893__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12894__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12894__A2 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12907__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12907__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12908__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12908__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12909__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12909__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12915__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12915__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12917__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12917__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12942__A1 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12943__A2 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12945__A1 (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12946__A1 (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12961__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12961__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12971__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12971__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12972__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12972__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12973__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12973__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12975__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12975__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12976__B (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12976__C (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12977__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12977__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12988__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12988__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12989__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12989__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12990__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12990__A2 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13003__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13003__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13004__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13004__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13005__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13005__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13011__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13011__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13012__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13012__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13013__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13013__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13026__A2 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13030__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13031__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13039__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13039__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13047__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13049__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13049__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13050__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13050__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13051__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13051__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13062__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13062__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13063__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13063__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13064__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13064__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13077__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13077__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13078__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13078__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13079__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13079__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13085__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13085__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13086__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13086__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13109__A1 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13114__A1 (.I(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13116__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13125__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13126__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13135__A1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13135__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13144__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13144__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13145__A1 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13145__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13156__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13156__A2 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13157__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13157__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13158__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13158__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13171__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13171__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13172__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13172__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13173__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13173__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13179__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13179__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13180__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13180__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13181__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13181__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13196__A2 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13203__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13206__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13207__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13212__A1 (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13217__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13217__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13237__A1 (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13237__A2 (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13237__A3 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13238__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13238__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13240__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13240__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13241__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13241__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13242__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13242__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13255__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13255__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13256__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13256__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13257__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13257__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13263__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13263__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13264__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13264__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13265__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13265__A2 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13284__A2 (.I(_06208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13286__A1 (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13287__A1 (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13287__B (.I(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13288__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13288__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13299__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13299__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13312__A1 (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13313__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13313__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13315__A1 (.I(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13315__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13317__A1 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13317__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13318__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13318__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13322__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13322__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13326__A1 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13334__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13334__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13335__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13335__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13344__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13344__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13345__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13345__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13346__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13346__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13360__A2 (.I(_06208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13364__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13365__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13365__A2 (.I(_06295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13366__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13369__A2 (.I(_06208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13386__A1 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13386__B (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13388__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13388__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13388__B (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13389__A1 (.I(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13389__A2 (.I(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13389__A3 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13391__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13391__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13395__A1 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13402__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13402__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13403__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13403__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13404__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13404__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13412__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13412__A2 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13413__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13413__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13414__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13414__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13433__A1 (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13436__A1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13437__A2 (.I(_06374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13451__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13451__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13456__A1 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13456__B (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13458__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13458__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13460__A1 (.I(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13460__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13466__A1 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13472__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13472__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13473__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13473__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13474__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13474__A2 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13482__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13482__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13483__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13483__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13484__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13484__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13496__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13500__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13501__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13501__A2 (.I(_06441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13507__B (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13508__A1 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13510__B2 (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13521__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13521__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13529__A1 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13529__B (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13533__A1 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13539__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13539__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13540__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13540__A2 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13541__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13541__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13547__A1 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13547__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13548__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13548__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13549__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13549__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13566__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13567__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13567__A2 (.I(_06512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13579__A1 (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13580__A1 (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13580__A2 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13586__A1 (.I(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13586__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13587__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13587__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13588__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13588__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13595__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13595__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13596__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13596__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13596__B (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13597__A1 (.I(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13597__A2 (.I(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13597__A3 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13608__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13608__A2 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13614__A2 (.I(_06563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13620__I0 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13620__I1 (.I(_06570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13620__S (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13622__A2 (.I(_06563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13629__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13629__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13635__A1 (.I(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13635__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13636__A1 (.I(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13636__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13646__A1 (.I(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13646__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13647__A1 (.I(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13647__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13653__A3 (.I(_06605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13658__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13658__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13659__A1 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13659__A2 (.I(_06611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13660__A1 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13660__A2 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13660__B (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13661__A1 (.I(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13661__A2 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13661__B (.I(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13662__A1 (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13662__A2 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13662__B (.I(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13663__A1 (.I(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13663__A2 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13663__B (.I(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13664__A1 (.I(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13664__A2 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13664__B (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13706__CLK (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13711__CLK (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13723__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13724__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13725__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13726__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13727__CLK (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13727__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13728__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13729__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13730__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13731__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13732__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13733__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13734__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13735__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13736__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13737__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13738__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13739__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13740__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13741__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13742__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13743__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13744__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13745__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13746__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13747__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13748__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13749__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13750__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13751__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13752__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13782__D (.I(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13784__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13785__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13786__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13787__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13788__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13789__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13790__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13791__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13792__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13793__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13794__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13795__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13796__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13797__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13798__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13799__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13800__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13801__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13803__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13804__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13805__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13806__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13807__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13808__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13809__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13810__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13811__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13812__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13813__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13814__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13815__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13816__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13817__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13848__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13849__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13850__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13851__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13852__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13853__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13854__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13855__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13856__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13857__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13858__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13859__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13860__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13861__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13862__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13863__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13864__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13865__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13866__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13867__CLK (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13867__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13868__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13869__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13870__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13871__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13872__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13873__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13874__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13875__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13876__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13877__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13878__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13879__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13880__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13881__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13882__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13883__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13884__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13885__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13886__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13887__CLK (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13887__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13888__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13889__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13890__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13891__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13892__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13893__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13894__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13895__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13896__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13897__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13898__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13899__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13900__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13901__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13902__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13903__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13904__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13905__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13906__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13907__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13908__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13909__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13910__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13911__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13912__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13913__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13914__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13915__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13916__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13917__CLK (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13917__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13918__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13919__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13920__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13921__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13922__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13923__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13924__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13925__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13926__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13927__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13928__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13929__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13930__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13931__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13932__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13933__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13934__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13935__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13936__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13937__CLK (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13937__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13938__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13939__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13940__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13941__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13942__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13943__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13944__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13945__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13946__CLK (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13946__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13947__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13948__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13949__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13950__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13951__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13952__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13953__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13954__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13955__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13956__RN (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13957__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone10_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone11_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone12_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone13_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone14_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone21_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone22_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone23_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone31_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone36_I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone39_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone43_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone44_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone48_I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone53_I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone54_I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone56_I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone57_I (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone59_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone6_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone7_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone8_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clone9_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout36_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold49_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold51_I (.I(FreqPhase[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold53_I (.I(FreqPhase[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold55_I (.I(FreqPhase[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold57_I (.I(FreqPhase[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold59_I (.I(FreqPhase[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold61_I (.I(FreqPhase[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold63_I (.I(FreqPhase[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold65_I (.I(FreqPhase[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold68_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold69_I (.I(FreqPhase[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold76_I (.I(LoadF));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold83_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold84_I (.I(FreqPhase[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold85_I (.I(FreqPhase[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold86_I (.I(FreqPhase[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold87_I (.I(FreqPhase[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold88_I (.I(FreqPhase[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold89_I (.I(FreqPhase[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold90_I (.I(LoadP));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold92_I (.I(Enable));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer25_I (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer32_I (.I(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer33_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer34_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer41_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer49_I (.I(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer62_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel DDS_Module_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_484 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06832_ (.I(\DDS_Stage.LCU.state[2] ),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06833_ (.A1(_05139_),
    .A2(\DDS_Stage.LCU.state[0] ),
    .A3(\DDS_Stage.LCU.state[1] ),
    .ZN(\DDS_Stage.LCU.SelMuxConfig ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06834_ (.A1(_05139_),
    .A2(\DDS_Stage.LCU.state[0] ),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 _06835_ (.I(net1),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 _06836_ (.I(_05171_),
    .Z(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06837_ (.I(net17),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06838_ (.A1(\DDS_Stage.LCU.state[2] ),
    .A2(\DDS_Stage.LCU.state[0] ),
    .A3(\DDS_Stage.LCU.state[1] ),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06839_ (.A1(_05182_),
    .A2(net18),
    .A3(_05193_),
    .A4(_05204_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06840_ (.I(\DDS_Stage.LCU.state[1] ),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06841_ (.A1(\DDS_Stage.LCU.state[2] ),
    .A2(\DDS_Stage.LCU.state[0] ),
    .A3(_05226_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06842_ (.A1(_05182_),
    .A2(net18),
    .A3(net17),
    .A4(_05237_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06843_ (.A1(\DDS_Stage.LCU.state[1] ),
    .A2(_05160_),
    .B(net125),
    .C(_05248_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06844_ (.I(_05171_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 _06845_ (.I(_05269_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06846_ (.A1(_05280_),
    .A2(net18),
    .A3(net17),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06847_ (.I(net18),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06848_ (.A1(_05280_),
    .A2(_05302_),
    .A3(_05193_),
    .B(_05237_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06849_ (.A1(\DDS_Stage.LCU.state[1] ),
    .A2(_05160_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06850_ (.A1(_05324_),
    .A2(_05291_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06851_ (.A1(_05182_),
    .A2(_05302_),
    .A3(net17),
    .A4(_05204_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06852_ (.A1(_05291_),
    .A2(_05313_),
    .B(_05335_),
    .C(net129),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06853_ (.A1(_05237_),
    .A2(net170),
    .Z(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06854_ (.I(_05366_),
    .Z(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 _06855_ (.I(_05171_),
    .Z(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06856_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-25] ),
    .Z(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 _06857_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[3] ),
    .Z(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 _06858_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[2] ),
    .Z(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _06859_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[0] ),
    .Z(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _06860_ (.I(_05431_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06861_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[1] ),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _06862_ (.I(_05452_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06863_ (.A1(_05442_),
    .A2(_05463_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06864_ (.A1(_05431_),
    .A2(_05452_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06865_ (.A1(_05474_),
    .A2(_05485_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06866_ (.A1(_05420_),
    .A2(_05496_),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06867_ (.A1(_05409_),
    .A2(_05507_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06868_ (.A1(_05420_),
    .A2(_05474_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06869_ (.A1(_05518_),
    .A2(_05529_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06870_ (.A1(_05431_),
    .A2(_05452_),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06871_ (.A1(_05420_),
    .A2(_05550_),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_16 _06872_ (.I(_05420_),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06873_ (.A1(_05572_),
    .A2(_05474_),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06874_ (.A1(_05561_),
    .A2(_05583_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06875_ (.A1(_05409_),
    .A2(_05594_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06876_ (.A1(_05171_),
    .A2(_05540_),
    .A3(_05605_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06877_ (.A1(_05387_),
    .A2(_05398_),
    .B(_05616_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06878_ (.I(_05627_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06879_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[4] ),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 _06880_ (.I(_05647_),
    .Z(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06881_ (.A1(_05442_),
    .A2(_05463_),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06882_ (.A1(_05550_),
    .A2(_05669_),
    .ZN(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06883_ (.A1(_05420_),
    .A2(_05680_),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06884_ (.A1(_05420_),
    .A2(_05463_),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06885_ (.A1(_05409_),
    .A2(_05702_),
    .ZN(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06886_ (.A1(_05691_),
    .A2(_05713_),
    .ZN(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06887_ (.A1(_05420_),
    .A2(_05474_),
    .ZN(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06888_ (.A1(_05409_),
    .A2(_05734_),
    .ZN(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06889_ (.A1(_05658_),
    .A2(_05724_),
    .A3(_05745_),
    .ZN(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06890_ (.A1(_05409_),
    .A2(_05529_),
    .B(_05658_),
    .ZN(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06891_ (.A1(_05572_),
    .A2(_05442_),
    .ZN(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06892_ (.A1(_05420_),
    .A2(_05485_),
    .ZN(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06893_ (.A1(_05767_),
    .A2(_05778_),
    .A3(_05789_),
    .ZN(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06894_ (.A1(_05387_),
    .A2(_05756_),
    .A3(_05800_),
    .ZN(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 _06895_ (.I(_05280_),
    .Z(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06896_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-24] ),
    .Z(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06897_ (.A1(_05822_),
    .A2(_05833_),
    .ZN(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06898_ (.A1(_05811_),
    .A2(_05844_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06899_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-23] ),
    .Z(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06900_ (.A1(_05420_),
    .A2(_05463_),
    .ZN(_05875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06901_ (.A1(_05431_),
    .A2(_05463_),
    .ZN(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06902_ (.A1(_05420_),
    .A2(_05886_),
    .ZN(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06903_ (.A1(_05572_),
    .A2(_05463_),
    .ZN(_05908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06904_ (.A1(_05897_),
    .A2(_05908_),
    .ZN(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06905_ (.A1(_05409_),
    .A2(_05919_),
    .ZN(_05930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06906_ (.A1(_05420_),
    .A2(_05431_),
    .ZN(_05940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06907_ (.A1(_05474_),
    .A2(_05940_),
    .ZN(_05951_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06908_ (.A1(_05409_),
    .A2(_05442_),
    .A3(_05875_),
    .B1(_05930_),
    .B2(_05951_),
    .ZN(_05962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06909_ (.A1(_05442_),
    .A2(_05452_),
    .ZN(_05973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06910_ (.A1(_05420_),
    .A2(_05973_),
    .ZN(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06911_ (.A1(_05420_),
    .A2(_05680_),
    .ZN(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06912_ (.A1(_05420_),
    .A2(_05886_),
    .B(_05995_),
    .C(_05409_),
    .ZN(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06913_ (.A1(_05409_),
    .A2(_05984_),
    .B(_06006_),
    .C(_05658_),
    .ZN(_06017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06914_ (.A1(_05658_),
    .A2(_05962_),
    .B(_06017_),
    .ZN(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06915_ (.I0(_05864_),
    .I1(_06028_),
    .S(_05182_),
    .Z(_06039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06916_ (.I(_06039_),
    .Z(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 _06917_ (.I(_05280_),
    .Z(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06918_ (.A1(_05442_),
    .A2(_05452_),
    .ZN(_06070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06919_ (.A1(_05420_),
    .A2(_06070_),
    .ZN(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06920_ (.A1(_05431_),
    .A2(_05463_),
    .ZN(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06921_ (.A1(_05409_),
    .A2(_06092_),
    .B(_05995_),
    .ZN(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06922_ (.A1(_05409_),
    .A2(_06081_),
    .B1(_06103_),
    .B2(_05529_),
    .ZN(_06114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06923_ (.A1(_05572_),
    .A2(_05442_),
    .ZN(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06924_ (.A1(_05658_),
    .A2(_06125_),
    .ZN(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_20 _06925_ (.I(_05647_),
    .ZN(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06926_ (.A1(_06146_),
    .A2(_06114_),
    .ZN(_06157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06927_ (.A1(_06114_),
    .A2(_06135_),
    .B(_06157_),
    .ZN(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06928_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-22] ),
    .Z(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06929_ (.A1(_05822_),
    .A2(_06179_),
    .ZN(_06190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06930_ (.A1(_06059_),
    .A2(_06168_),
    .B(_06190_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06931_ (.A1(_05420_),
    .A2(_05442_),
    .ZN(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06932_ (.A1(_05409_),
    .A2(_06211_),
    .ZN(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_16 _06933_ (.I(_05409_),
    .ZN(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06934_ (.A1(_05572_),
    .A2(_05886_),
    .ZN(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06935_ (.A1(_06232_),
    .A2(_05875_),
    .A3(_06243_),
    .ZN(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06936_ (.A1(_05734_),
    .A2(_06221_),
    .B(_06254_),
    .ZN(_06265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06937_ (.A1(_06146_),
    .A2(_05529_),
    .ZN(_06276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06938_ (.A1(_05658_),
    .A2(_06265_),
    .ZN(_06287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06939_ (.A1(_06265_),
    .A2(_06276_),
    .B(_06287_),
    .ZN(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06940_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-21] ),
    .Z(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06941_ (.A1(_05822_),
    .A2(_06308_),
    .ZN(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06942_ (.A1(_06059_),
    .A2(_06297_),
    .B(_06319_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06943_ (.A1(_05420_),
    .A2(_05496_),
    .ZN(_06340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06944_ (.A1(_05583_),
    .A2(_06340_),
    .ZN(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06945_ (.A1(_05409_),
    .A2(_06351_),
    .ZN(_06362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06946_ (.A1(_05420_),
    .A2(_05496_),
    .B(_05409_),
    .ZN(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06947_ (.A1(_05778_),
    .A2(_06373_),
    .ZN(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06948_ (.A1(_06362_),
    .A2(_06383_),
    .ZN(_06394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06949_ (.A1(_06146_),
    .A2(_06394_),
    .Z(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06950_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-20] ),
    .Z(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06951_ (.A1(_05822_),
    .A2(net152),
    .ZN(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06952_ (.A1(_06059_),
    .A2(_06405_),
    .B(_06427_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06953_ (.A1(_05572_),
    .A2(_05680_),
    .ZN(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06954_ (.A1(_05572_),
    .A2(_05463_),
    .ZN(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06955_ (.A1(_05409_),
    .A2(_06458_),
    .ZN(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06956_ (.I(_05691_),
    .ZN(_06480_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06957_ (.A1(_06232_),
    .A2(_06480_),
    .A3(_06081_),
    .ZN(_06491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06958_ (.A1(_06447_),
    .A2(_06469_),
    .B(_06491_),
    .ZN(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06959_ (.A1(_06146_),
    .A2(_06502_),
    .Z(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06960_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-19] ),
    .Z(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06961_ (.A1(_05822_),
    .A2(net155),
    .ZN(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06962_ (.A1(_06059_),
    .A2(_06513_),
    .B(_06534_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06963_ (.A1(_05572_),
    .A2(_06092_),
    .ZN(_06555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06964_ (.A1(_05409_),
    .A2(_05908_),
    .ZN(_06566_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _06965_ (.A1(_05409_),
    .A2(_06081_),
    .A3(_06555_),
    .B1(_06566_),
    .B2(_05431_),
    .ZN(_06576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06966_ (.A1(_05658_),
    .A2(_06576_),
    .Z(_06587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06967_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-18] ),
    .Z(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06968_ (.A1(_05822_),
    .A2(_06598_),
    .ZN(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06969_ (.A1(_06059_),
    .A2(_06587_),
    .B(_06609_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06970_ (.A1(_05409_),
    .A2(_05951_),
    .ZN(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06971_ (.A1(_05550_),
    .A2(_05778_),
    .ZN(_06614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06972_ (.A1(_05713_),
    .A2(_06614_),
    .ZN(_06615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06973_ (.A1(_05919_),
    .A2(_06613_),
    .B(_06615_),
    .ZN(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06974_ (.A1(_05658_),
    .A2(_06616_),
    .Z(_06617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06975_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-17] ),
    .Z(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06976_ (.A1(_05822_),
    .A2(_06618_),
    .ZN(_06619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06977_ (.A1(_06059_),
    .A2(_06617_),
    .B(_06619_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06978_ (.I(_05908_),
    .ZN(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06979_ (.A1(_05420_),
    .A2(_05431_),
    .ZN(_06621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06980_ (.A1(_05409_),
    .A2(_06621_),
    .ZN(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06981_ (.A1(_05420_),
    .A2(_05973_),
    .ZN(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06982_ (.A1(_06232_),
    .A2(_06620_),
    .ZN(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06983_ (.A1(_06620_),
    .A2(_06622_),
    .B(_06623_),
    .C(_06624_),
    .ZN(_06625_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06984_ (.A1(_06146_),
    .A2(_06625_),
    .Z(_06626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06985_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-16] ),
    .Z(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06986_ (.A1(_05822_),
    .A2(_06627_),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06987_ (.A1(_06059_),
    .A2(_06626_),
    .B(_06628_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06988_ (.A1(_05409_),
    .A2(_05778_),
    .ZN(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06989_ (.A1(_05583_),
    .A2(_06469_),
    .ZN(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06990_ (.A1(_06629_),
    .A2(_06630_),
    .ZN(_06631_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06991_ (.A1(_05658_),
    .A2(_06631_),
    .Z(_06632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06992_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-15] ),
    .Z(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06993_ (.A1(_05822_),
    .A2(_06633_),
    .ZN(_06634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06994_ (.A1(_06059_),
    .A2(_06632_),
    .B(_06634_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06995_ (.A1(_05507_),
    .A2(_06221_),
    .B(_06383_),
    .ZN(_06635_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06996_ (.A1(_06146_),
    .A2(_06635_),
    .Z(_06636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _06997_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-14] ),
    .Z(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06998_ (.A1(_05822_),
    .A2(_06637_),
    .ZN(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06999_ (.A1(_06059_),
    .A2(_06636_),
    .B(_06638_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07000_ (.A1(_05409_),
    .A2(_05572_),
    .ZN(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07001_ (.A1(_05647_),
    .A2(_05485_),
    .Z(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07002_ (.A1(_06639_),
    .A2(_06640_),
    .Z(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _07003_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-13] ),
    .Z(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07004_ (.A1(_05822_),
    .A2(_06642_),
    .ZN(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07005_ (.A1(_06059_),
    .A2(_06641_),
    .B(_06643_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07006_ (.A1(_06243_),
    .A2(_06623_),
    .ZN(_06644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07007_ (.A1(_05420_),
    .A2(_05452_),
    .ZN(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07008_ (.A1(_05409_),
    .A2(_05431_),
    .A3(_06645_),
    .ZN(_06646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07009_ (.A1(_05409_),
    .A2(_06644_),
    .B(_06646_),
    .ZN(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07010_ (.A1(_06146_),
    .A2(_06647_),
    .Z(_06648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07011_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-12] ),
    .Z(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07012_ (.A1(_05822_),
    .A2(_06649_),
    .ZN(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07013_ (.A1(_06059_),
    .A2(_06648_),
    .B(_06650_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07014_ (.A1(_05572_),
    .A2(_05452_),
    .ZN(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07015_ (.A1(_06651_),
    .A2(_06629_),
    .ZN(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07016_ (.A1(_06146_),
    .A2(_06652_),
    .Z(_06653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07017_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-11] ),
    .Z(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07018_ (.A1(_05822_),
    .A2(_06654_),
    .ZN(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07019_ (.A1(_06059_),
    .A2(_06653_),
    .B(_06655_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07020_ (.A1(_05409_),
    .A2(_05940_),
    .ZN(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07021_ (.A1(_06615_),
    .A2(_06656_),
    .ZN(_06657_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07022_ (.A1(_05658_),
    .A2(_06657_),
    .Z(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _07023_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-10] ),
    .Z(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07024_ (.A1(_05822_),
    .A2(_06659_),
    .ZN(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07025_ (.A1(_06059_),
    .A2(_06658_),
    .B(_06660_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07026_ (.A1(_05409_),
    .A2(_05420_),
    .A3(_05474_),
    .ZN(_06661_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07027_ (.A1(_05583_),
    .A2(_06211_),
    .A3(_06661_),
    .ZN(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07028_ (.A1(_06146_),
    .A2(_06662_),
    .Z(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07029_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-9] ),
    .Z(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07030_ (.A1(_05822_),
    .A2(_06664_),
    .ZN(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07031_ (.A1(_06059_),
    .A2(_06663_),
    .B(_06665_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07032_ (.A1(_05572_),
    .A2(_05669_),
    .ZN(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07033_ (.A1(_05897_),
    .A2(_06666_),
    .ZN(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07034_ (.A1(_05647_),
    .A2(_05409_),
    .Z(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07035_ (.A1(_05680_),
    .A2(_06668_),
    .ZN(_06669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07036_ (.A1(_05658_),
    .A2(_05680_),
    .B(_06669_),
    .ZN(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07037_ (.A1(_06667_),
    .A2(_06670_),
    .Z(_06671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _07038_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-8] ),
    .Z(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07039_ (.A1(_05822_),
    .A2(_06672_),
    .ZN(_06673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07040_ (.A1(_06059_),
    .A2(_06671_),
    .B(_06673_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07041_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-7] ),
    .Z(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07042_ (.A1(_05822_),
    .A2(_06674_),
    .ZN(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07043_ (.A1(_06059_),
    .A2(_06640_),
    .B(_06675_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07044_ (.A1(_05518_),
    .A2(_06340_),
    .ZN(_06676_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07045_ (.A1(_06232_),
    .A2(_05702_),
    .A3(_06555_),
    .B(_06676_),
    .ZN(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07046_ (.A1(_05658_),
    .A2(_06677_),
    .Z(_06678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07047_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-6] ),
    .Z(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07048_ (.A1(_05822_),
    .A2(_06679_),
    .ZN(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07049_ (.A1(_06059_),
    .A2(_06678_),
    .B(_06680_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07050_ (.A1(_06232_),
    .A2(_05485_),
    .ZN(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07051_ (.A1(_05583_),
    .A2(_06681_),
    .ZN(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07052_ (.A1(_06624_),
    .A2(_06682_),
    .ZN(_06683_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07053_ (.A1(_06146_),
    .A2(_06683_),
    .Z(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07054_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-5] ),
    .Z(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07055_ (.A1(_05822_),
    .A2(_06685_),
    .ZN(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07056_ (.A1(_06059_),
    .A2(_06684_),
    .B(_06686_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07057_ (.A1(_06232_),
    .A2(_06620_),
    .ZN(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07058_ (.A1(_05409_),
    .A2(_06125_),
    .ZN(_06688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07059_ (.A1(_06687_),
    .A2(_06688_),
    .ZN(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07060_ (.A1(_05658_),
    .A2(_06689_),
    .Z(_06690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07061_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-4] ),
    .Z(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07062_ (.A1(_05822_),
    .A2(_06691_),
    .ZN(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07063_ (.A1(_06059_),
    .A2(_06690_),
    .B(_06692_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07064_ (.A1(_05420_),
    .A2(_06681_),
    .ZN(_06693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07065_ (.A1(_05409_),
    .A2(_05594_),
    .B(_06693_),
    .ZN(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07066_ (.A1(_05658_),
    .A2(_06694_),
    .Z(_06695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07067_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-3] ),
    .Z(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07068_ (.A1(_05822_),
    .A2(_06696_),
    .ZN(_06697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07069_ (.A1(_06059_),
    .A2(_06695_),
    .B(_06697_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07070_ (.A1(_05409_),
    .A2(_06340_),
    .ZN(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07071_ (.A1(_05409_),
    .A2(_05485_),
    .B1(_05507_),
    .B2(_06698_),
    .ZN(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07072_ (.A1(_05658_),
    .A2(_06699_),
    .Z(_06700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07073_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-2] ),
    .Z(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07074_ (.A1(_05822_),
    .A2(_06701_),
    .ZN(_06702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07075_ (.A1(_06059_),
    .A2(_06700_),
    .B(_06702_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07076_ (.A1(_05572_),
    .A2(_05452_),
    .ZN(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07077_ (.A1(_05409_),
    .A2(_06651_),
    .ZN(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07078_ (.A1(_06703_),
    .A2(_06704_),
    .ZN(_06705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07079_ (.A1(_05930_),
    .A2(_06705_),
    .ZN(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07080_ (.A1(_05658_),
    .A2(_06706_),
    .Z(_06707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07081_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-1] ),
    .Z(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07082_ (.A1(_05822_),
    .A2(_06708_),
    .ZN(_06709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07083_ (.A1(_06059_),
    .A2(_06707_),
    .B(_06709_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07084_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[0] ),
    .Z(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07085_ (.A1(_05420_),
    .A2(_05669_),
    .B(_05409_),
    .ZN(_06711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07086_ (.A1(_06243_),
    .A2(_06711_),
    .ZN(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07087_ (.A1(_05572_),
    .A2(_05550_),
    .ZN(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07088_ (.A1(_05420_),
    .A2(_06070_),
    .ZN(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07089_ (.A1(_06713_),
    .A2(_06714_),
    .ZN(_06715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07090_ (.A1(_05409_),
    .A2(_06715_),
    .ZN(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07091_ (.A1(_06712_),
    .A2(_06716_),
    .ZN(_06717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07092_ (.A1(_05658_),
    .A2(_06717_),
    .Z(_06718_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07093_ (.I0(_06710_),
    .I1(_06718_),
    .S(_05182_),
    .Z(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07094_ (.I(_06719_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07095_ (.A1(_05420_),
    .A2(_06092_),
    .ZN(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07096_ (.A1(_05420_),
    .A2(_05886_),
    .B(_06232_),
    .ZN(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07097_ (.A1(_06720_),
    .A2(_06721_),
    .ZN(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07098_ (.A1(_06146_),
    .A2(_06722_),
    .Z(_06723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07099_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[1] ),
    .Z(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07100_ (.A1(_05822_),
    .A2(_06724_),
    .ZN(_06725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07101_ (.A1(_06059_),
    .A2(_06723_),
    .B(_06725_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07102_ (.A1(_05572_),
    .A2(_05431_),
    .ZN(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07103_ (.A1(_05420_),
    .A2(_05485_),
    .B(_06232_),
    .ZN(_06727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07104_ (.A1(_06713_),
    .A2(_06688_),
    .B1(_06726_),
    .B2(_06727_),
    .ZN(_06728_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07105_ (.A1(_06146_),
    .A2(_06728_),
    .Z(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07106_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[2] ),
    .Z(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07107_ (.A1(_05822_),
    .A2(_06730_),
    .ZN(_06731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07108_ (.A1(_06059_),
    .A2(_06729_),
    .B(_06731_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07109_ (.A1(_06713_),
    .A2(_06645_),
    .ZN(_06732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07110_ (.A1(_05420_),
    .A2(_05669_),
    .ZN(_06733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07111_ (.A1(_05908_),
    .A2(_06733_),
    .ZN(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07112_ (.A1(_05409_),
    .A2(_06734_),
    .ZN(_06735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07113_ (.A1(_05409_),
    .A2(_06732_),
    .B(_06735_),
    .ZN(_06736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07114_ (.A1(_05658_),
    .A2(_06736_),
    .Z(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07115_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[3] ),
    .Z(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07116_ (.A1(_05822_),
    .A2(_06738_),
    .ZN(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07117_ (.A1(_06059_),
    .A2(_06737_),
    .B(_06739_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07118_ (.A1(_06092_),
    .A2(_06622_),
    .B(_06713_),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07119_ (.A1(_05658_),
    .A2(_06740_),
    .Z(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _07120_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[4] ),
    .Z(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07121_ (.A1(_05822_),
    .A2(_06742_),
    .ZN(_06743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07122_ (.A1(_06059_),
    .A2(_06741_),
    .B(_06743_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07123_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[5] ),
    .Z(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07124_ (.A1(_05280_),
    .A2(_06744_),
    .ZN(_06745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07125_ (.A1(_06059_),
    .A2(_06668_),
    .B(_06745_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07126_ (.A1(_05409_),
    .A2(_05778_),
    .A3(_05789_),
    .ZN(_06746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07127_ (.A1(_05658_),
    .A2(_05540_),
    .A3(_06746_),
    .ZN(_06747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07128_ (.A1(_05572_),
    .A2(_05431_),
    .B(_05409_),
    .ZN(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07129_ (.A1(_05897_),
    .A2(_06748_),
    .ZN(_06749_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07130_ (.A1(_05431_),
    .A2(_06566_),
    .B(_06749_),
    .C(_06146_),
    .ZN(_06750_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07131_ (.A1(_05387_),
    .A2(_06747_),
    .A3(_06750_),
    .ZN(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07132_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-25] ),
    .ZN(_06752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07133_ (.A1(_06751_),
    .A2(_06752_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07134_ (.A1(_05572_),
    .A2(_06092_),
    .ZN(_06753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07135_ (.A1(_06232_),
    .A2(_06458_),
    .ZN(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07136_ (.A1(_06753_),
    .A2(_06754_),
    .ZN(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07137_ (.A1(_05572_),
    .A2(_05485_),
    .ZN(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07138_ (.A1(_06469_),
    .A2(_06756_),
    .ZN(_06757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07139_ (.A1(_06755_),
    .A2(_06757_),
    .B(_05658_),
    .ZN(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07140_ (.A1(_06232_),
    .A2(_05463_),
    .ZN(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07141_ (.A1(_05431_),
    .A2(_06759_),
    .B(_05420_),
    .ZN(_06760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07142_ (.A1(_05409_),
    .A2(_05452_),
    .ZN(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07143_ (.A1(_05658_),
    .A2(_06761_),
    .ZN(_06762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07144_ (.A1(_06760_),
    .A2(_06762_),
    .B(_05171_),
    .ZN(_06763_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07145_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-24] ),
    .B1(_06758_),
    .B2(_06763_),
    .ZN(_06764_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07146_ (.I(_06764_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07147_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-23] ),
    .ZN(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07148_ (.A1(_06447_),
    .A2(_06688_),
    .ZN(_06766_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07149_ (.A1(_06146_),
    .A2(_06716_),
    .A3(_06766_),
    .Z(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07150_ (.A1(_06243_),
    .A2(_06469_),
    .B(_06146_),
    .ZN(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07151_ (.A1(_06232_),
    .A2(_06734_),
    .B(_06768_),
    .ZN(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07152_ (.A1(_05182_),
    .A2(_06769_),
    .ZN(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07153_ (.A1(_05387_),
    .A2(_06765_),
    .B1(_06767_),
    .B2(_06770_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07154_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-22] ),
    .ZN(_06771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07155_ (.A1(_05409_),
    .A2(_06732_),
    .ZN(_06772_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07156_ (.A1(_05658_),
    .A2(_06766_),
    .A3(_06772_),
    .ZN(_06773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07157_ (.A1(_05409_),
    .A2(_06726_),
    .ZN(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07158_ (.A1(_06092_),
    .A2(_06774_),
    .B(_06757_),
    .C(_06146_),
    .ZN(_06775_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07159_ (.A1(_05387_),
    .A2(_06773_),
    .A3(_06775_),
    .ZN(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07160_ (.A1(_06771_),
    .A2(_06776_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07161_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-21] ),
    .ZN(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07162_ (.A1(_05409_),
    .A2(_05789_),
    .ZN(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07163_ (.A1(_05409_),
    .A2(_06651_),
    .A3(_05875_),
    .ZN(_06779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07164_ (.A1(_06232_),
    .A2(_06644_),
    .B(_05658_),
    .ZN(_06780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07165_ (.A1(_05431_),
    .A2(_06779_),
    .B(_06780_),
    .ZN(_06781_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07166_ (.A1(_06146_),
    .A2(_06778_),
    .B(_06781_),
    .C(_05182_),
    .ZN(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07167_ (.A1(_05387_),
    .A2(_06777_),
    .B(_06782_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07168_ (.A1(_05724_),
    .A2(_06629_),
    .B(_06146_),
    .ZN(_06783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07169_ (.A1(_05550_),
    .A2(_06681_),
    .B(_06373_),
    .C(_05658_),
    .ZN(_06784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07170_ (.A1(_06783_),
    .A2(_06784_),
    .B(_05182_),
    .ZN(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07171_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-20] ),
    .ZN(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07172_ (.A1(_06785_),
    .A2(_06786_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07173_ (.A1(_05420_),
    .A2(_05886_),
    .ZN(_06787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07174_ (.A1(_05409_),
    .A2(_05875_),
    .ZN(_06788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07175_ (.A1(_05420_),
    .A2(_05485_),
    .B(_05409_),
    .ZN(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07176_ (.A1(_06726_),
    .A2(_06789_),
    .ZN(_06790_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07177_ (.A1(_06787_),
    .A2(_06788_),
    .B(_05658_),
    .C(_06790_),
    .ZN(_06791_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07178_ (.A1(_06146_),
    .A2(_05886_),
    .A3(_06645_),
    .A4(_06629_),
    .ZN(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07179_ (.A1(_05182_),
    .A2(_06791_),
    .A3(_06792_),
    .ZN(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07180_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-19] ),
    .ZN(_06794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07181_ (.A1(_06793_),
    .A2(_06794_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07182_ (.A1(_05409_),
    .A2(_05529_),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07183_ (.A1(_05507_),
    .A2(_06795_),
    .B(_05647_),
    .ZN(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07184_ (.I(_06796_),
    .ZN(_06797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07185_ (.A1(_05452_),
    .A2(_06748_),
    .ZN(_06798_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07186_ (.A1(_05409_),
    .A2(_06651_),
    .A3(_06340_),
    .ZN(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07187_ (.A1(_06797_),
    .A2(_06798_),
    .B1(_06799_),
    .B2(_06780_),
    .ZN(_06800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07188_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-18] ),
    .I1(_06800_),
    .S(_05182_),
    .Z(_06801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07189_ (.I(_06801_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07190_ (.A1(_05409_),
    .A2(_05550_),
    .B(_05691_),
    .ZN(_06802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07191_ (.A1(_05658_),
    .A2(_06681_),
    .ZN(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07192_ (.A1(_05658_),
    .A2(_06802_),
    .B1(_06803_),
    .B2(_06715_),
    .ZN(_06804_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07193_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-17] ),
    .I1(_06804_),
    .S(_05182_),
    .Z(_06805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07194_ (.I(_06805_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07195_ (.A1(_05409_),
    .A2(_05452_),
    .ZN(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07196_ (.A1(_05702_),
    .A2(_06806_),
    .B(_05658_),
    .C(_05669_),
    .ZN(_06807_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07197_ (.A1(_06726_),
    .A2(_06759_),
    .B1(_06774_),
    .B2(_06703_),
    .C(_06146_),
    .ZN(_06808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07198_ (.A1(_06807_),
    .A2(_06808_),
    .ZN(_06809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07199_ (.A1(_05182_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-16] ),
    .ZN(_06810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07200_ (.A1(_05387_),
    .A2(_06809_),
    .B(_06810_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07201_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-15] ),
    .ZN(_06811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07202_ (.A1(_05518_),
    .A2(_06340_),
    .B1(_06721_),
    .B2(_05778_),
    .C(_05658_),
    .ZN(_06812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07203_ (.A1(_05420_),
    .A2(_05550_),
    .B(_06774_),
    .ZN(_06813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07204_ (.A1(_06646_),
    .A2(_06813_),
    .B(_05658_),
    .ZN(_06814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07205_ (.A1(_05182_),
    .A2(_06814_),
    .ZN(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07206_ (.A1(_05387_),
    .A2(_06811_),
    .B1(_06812_),
    .B2(_06815_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07207_ (.A1(_06232_),
    .A2(_05431_),
    .B(_05658_),
    .ZN(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07208_ (.A1(_06362_),
    .A2(_06768_),
    .B1(_06816_),
    .B2(_06761_),
    .ZN(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07209_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-14] ),
    .I1(_06817_),
    .S(_05182_),
    .Z(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07210_ (.I(_06818_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07211_ (.A1(_05409_),
    .A2(_06555_),
    .A3(_06787_),
    .ZN(_06819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07212_ (.A1(_05658_),
    .A2(_06755_),
    .ZN(_06820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07213_ (.A1(_06713_),
    .A2(_06681_),
    .B1(_06748_),
    .B2(_05496_),
    .ZN(_06821_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _07214_ (.A1(_06819_),
    .A2(_06820_),
    .B1(_06821_),
    .B2(_05658_),
    .C(_05171_),
    .ZN(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07215_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-13] ),
    .B(_06822_),
    .ZN(_06823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07216_ (.I(_06823_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07217_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-12] ),
    .ZN(_06824_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07218_ (.A1(_05409_),
    .A2(_05550_),
    .B1(_06092_),
    .B2(_06622_),
    .C(_05658_),
    .ZN(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07219_ (.A1(_05669_),
    .A2(_06688_),
    .ZN(_06826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07220_ (.A1(_05409_),
    .A2(_06614_),
    .B(_05658_),
    .ZN(_06827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07221_ (.A1(_06826_),
    .A2(_06827_),
    .ZN(_06828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07222_ (.A1(_05182_),
    .A2(_06825_),
    .A3(_06828_),
    .ZN(_06829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07223_ (.A1(_05387_),
    .A2(_06824_),
    .B(_06829_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07224_ (.A1(_05409_),
    .A2(_05485_),
    .A3(_05594_),
    .ZN(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07225_ (.A1(_06232_),
    .A2(_06211_),
    .A3(_06756_),
    .Z(_06831_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _07226_ (.A1(_05658_),
    .A2(_06681_),
    .A3(_06830_),
    .B1(_06831_),
    .B2(_06796_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07227_ (.A1(_05182_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-11] ),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07228_ (.A1(_05387_),
    .A2(_00292_),
    .B(_00293_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07229_ (.A1(_06714_),
    .A2(_06666_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07230_ (.A1(_05409_),
    .A2(_00294_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07231_ (.A1(_05658_),
    .A2(_06125_),
    .B(_06749_),
    .C(_00295_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07232_ (.A1(_05182_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-10] ),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07233_ (.A1(_05387_),
    .A2(_00296_),
    .B(_00297_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07234_ (.A1(_06211_),
    .A2(_06687_),
    .B(_06146_),
    .C(_06006_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07235_ (.A1(_05409_),
    .A2(_06211_),
    .A3(_06756_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07236_ (.A1(_06624_),
    .A2(_00299_),
    .B(_05658_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07237_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-9] ),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07238_ (.A1(_05822_),
    .A2(_00298_),
    .A3(_00300_),
    .B(_00301_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07239_ (.A1(_06651_),
    .A2(_06714_),
    .B(_05409_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07240_ (.A1(_05658_),
    .A2(_06698_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _07241_ (.A1(_05409_),
    .A2(_06720_),
    .B1(_06774_),
    .B2(_06480_),
    .C(_06146_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07242_ (.A1(_00302_),
    .A2(_00303_),
    .B(_00304_),
    .C(_05182_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07243_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-8] ),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07244_ (.A1(_00305_),
    .A2(_00306_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07245_ (.A1(_05518_),
    .A2(_06211_),
    .B1(_06732_),
    .B2(_05409_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07246_ (.A1(_06232_),
    .A2(_05474_),
    .B(_05658_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07247_ (.A1(_05409_),
    .A2(_06447_),
    .A3(_06733_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07248_ (.A1(_05658_),
    .A2(_00307_),
    .B1(_00308_),
    .B2(_00309_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07249_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-7] ),
    .I1(_00310_),
    .S(_05182_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07250_ (.I(_00311_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07251_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-6] ),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07252_ (.A1(_06232_),
    .A2(_06351_),
    .B1(_06681_),
    .B2(_05550_),
    .C(_05658_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07253_ (.A1(_05658_),
    .A2(_06623_),
    .A3(_06735_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07254_ (.A1(_05182_),
    .A2(_00314_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07255_ (.A1(_05387_),
    .A2(_00312_),
    .B1(_00313_),
    .B2(_00315_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07256_ (.A1(_05431_),
    .A2(_05713_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07257_ (.A1(_05658_),
    .A2(_00316_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07258_ (.A1(_06146_),
    .A2(_06623_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07259_ (.A1(_06491_),
    .A2(_00317_),
    .B1(_00318_),
    .B2(_06629_),
    .C(_05171_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07260_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-5] ),
    .B(_00319_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07261_ (.I(_00320_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07262_ (.A1(_05409_),
    .A2(_05691_),
    .B(_05767_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07263_ (.A1(_05409_),
    .A2(_05875_),
    .A3(_06666_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07264_ (.A1(_05658_),
    .A2(_06826_),
    .A3(_00322_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07265_ (.A1(_00321_),
    .A2(_00323_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07266_ (.A1(_05182_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-4] ),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07267_ (.A1(_05387_),
    .A2(_00324_),
    .B(_00325_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07268_ (.A1(_06232_),
    .A2(_06125_),
    .B1(_06727_),
    .B2(_06753_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07269_ (.A1(_05409_),
    .A2(_05485_),
    .A3(_05561_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _07270_ (.A1(_05658_),
    .A2(_00326_),
    .B1(_00327_),
    .B2(_06762_),
    .C(_05171_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07271_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-3] ),
    .B(_00328_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07272_ (.I(_00329_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07273_ (.A1(_05409_),
    .A2(_05431_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07274_ (.A1(_06651_),
    .A2(_00330_),
    .B1(_06759_),
    .B2(_05431_),
    .C(_06146_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07275_ (.A1(_06232_),
    .A2(_06645_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07276_ (.A1(_05995_),
    .A2(_06622_),
    .B(_00332_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07277_ (.A1(_06146_),
    .A2(_00333_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07278_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-2] ),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07279_ (.A1(_05822_),
    .A2(_00331_),
    .A3(_00334_),
    .B(_00335_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07280_ (.A1(_05734_),
    .A2(_06681_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07281_ (.A1(_05658_),
    .A2(_06624_),
    .A3(_00336_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07282_ (.A1(_06081_),
    .A2(_06788_),
    .B(_06146_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07283_ (.A1(_05182_),
    .A2(_00337_),
    .A3(_00338_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07284_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-1] ),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07285_ (.A1(_00339_),
    .A2(_00340_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07286_ (.A1(_05583_),
    .A2(_06711_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07287_ (.A1(_00295_),
    .A2(_00341_),
    .B(_06146_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07288_ (.A1(_05409_),
    .A2(_05702_),
    .B(_05658_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07289_ (.A1(_00342_),
    .A2(_00343_),
    .B(_05182_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07290_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[0] ),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07291_ (.A1(_00344_),
    .A2(_00345_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07292_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[1] ),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07293_ (.A1(_05409_),
    .A2(_06555_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07294_ (.A1(_05658_),
    .A2(_06232_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07295_ (.A1(_06491_),
    .A2(_00347_),
    .A3(_00348_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07296_ (.A1(_05658_),
    .A2(_06687_),
    .B(_05171_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07297_ (.A1(_05387_),
    .A2(_00346_),
    .B1(_00349_),
    .B2(_00350_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07298_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-15] ),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07299_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-15] ),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07300_ (.I0(net66),
    .I1(net58),
    .S(_05182_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07301_ (.I(_00353_),
    .Z(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07302_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-14] ),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 _07303_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-14] ),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07304_ (.I0(net54),
    .I1(_00355_),
    .S(_05182_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07305_ (.I(_00356_),
    .Z(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07306_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-13] ),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _07307_ (.I(net161),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07308_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-13] ),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07309_ (.A1(_05280_),
    .A2(net70),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07310_ (.A1(_06059_),
    .A2(_00358_),
    .B(_00360_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 _07311_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-12] ),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07312_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-12] ),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 _07313_ (.I(_00362_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07314_ (.I0(_00361_),
    .I1(net60),
    .S(_05182_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07315_ (.I(_00364_),
    .Z(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 _07316_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-11] ),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07317_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-11] ),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07318_ (.I(_00366_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07319_ (.I0(_00365_),
    .I1(net61),
    .S(_05182_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07320_ (.I(_00368_),
    .Z(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07321_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-10] ),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07322_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-10] ),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07323_ (.I0(_00369_),
    .I1(_00370_),
    .S(_05182_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07324_ (.I(_00371_),
    .Z(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 _07325_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-9] ),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 _07326_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-9] ),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07327_ (.I0(_00372_),
    .I1(_00373_),
    .S(_05182_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07328_ (.I(_00374_),
    .Z(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07329_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-8] ),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07330_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-8] ),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07331_ (.I0(_00375_),
    .I1(_00376_),
    .S(_05182_),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07332_ (.I(_00377_),
    .Z(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07333_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-7] ),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07334_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-7] ),
    .Z(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07335_ (.I0(_00378_),
    .I1(_00379_),
    .S(_05182_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07336_ (.I(_00380_),
    .Z(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 _07337_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-6] ),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 _07338_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-6] ),
    .Z(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07339_ (.I0(_00381_),
    .I1(_00382_),
    .S(_05182_),
    .Z(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07340_ (.I(_00383_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 _07341_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-5] ),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 _07342_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-5] ),
    .Z(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07343_ (.I0(_00384_),
    .I1(_00385_),
    .S(_05182_),
    .Z(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07344_ (.I(_00386_),
    .Z(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07345_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-4] ),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07346_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-4] ),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07347_ (.I0(_00387_),
    .I1(_00388_),
    .S(_05182_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07348_ (.I(_00389_),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07349_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-3] ),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 _07350_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-3] ),
    .Z(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07351_ (.I0(_00390_),
    .I1(net63),
    .S(_05182_),
    .Z(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07352_ (.I(_00392_),
    .Z(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 _07353_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-2] ),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 _07354_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-2] ),
    .Z(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 _07355_ (.I(_05171_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07356_ (.I0(_00393_),
    .I1(_00394_),
    .S(_00395_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07357_ (.I(_00396_),
    .Z(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 _07358_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-1] ),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 _07359_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-1] ),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07360_ (.I0(_00397_),
    .I1(_00398_),
    .S(_00395_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07361_ (.I(_00399_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07362_ (.A1(\DDS_Stage.LCU.state[2] ),
    .A2(_05226_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07363_ (.A1(\DDS_Stage.LCU.state[0] ),
    .A2(_00400_),
    .B(\DDS_Stage.LCU.SelMuxConfig ),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 _07364_ (.I(_00401_),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07365_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-15] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-15] ),
    .S(_00402_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07366_ (.I(_00403_),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07367_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-14] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-14] ),
    .S(_00402_),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07368_ (.I(_00404_),
    .Z(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07369_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-13] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-13] ),
    .S(_00402_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07370_ (.I(_00405_),
    .Z(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07371_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-12] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-12] ),
    .S(_00402_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07372_ (.I(_00406_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07373_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-11] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-11] ),
    .S(_00402_),
    .Z(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07374_ (.I(_00407_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07375_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-10] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-10] ),
    .S(_00402_),
    .Z(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07376_ (.I(_00408_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07377_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-9] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-9] ),
    .S(_00402_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07378_ (.I(_00409_),
    .Z(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07379_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-8] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-8] ),
    .S(_00402_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07380_ (.I(_00410_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07381_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-7] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-7] ),
    .S(_00402_),
    .Z(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07382_ (.I(_00411_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07383_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-6] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-6] ),
    .S(_00402_),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07384_ (.I(_00412_),
    .Z(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07385_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-5] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-5] ),
    .S(_00402_),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07386_ (.I(_00413_),
    .Z(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07387_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-4] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-4] ),
    .S(_00402_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07388_ (.I(_00414_),
    .Z(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07389_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-3] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-3] ),
    .S(_00402_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07390_ (.I(_00415_),
    .Z(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07391_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-2] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-2] ),
    .S(_00402_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07392_ (.I(_00416_),
    .Z(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07393_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-1] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-1] ),
    .S(_00402_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07394_ (.I(_00417_),
    .Z(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07395_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-25] ),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07396_ (.A1(_05409_),
    .A2(_06714_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07397_ (.A1(_05658_),
    .A2(_06779_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07398_ (.A1(_05409_),
    .A2(_05897_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07399_ (.A1(_05995_),
    .A2(_00421_),
    .B(_06254_),
    .C(_06146_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07400_ (.A1(_00419_),
    .A2(_00420_),
    .B(_00422_),
    .C(_05182_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07401_ (.A1(_05387_),
    .A2(_00418_),
    .B(_00423_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07402_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-24] ),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07403_ (.A1(_05529_),
    .A2(_06666_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07404_ (.A1(_06668_),
    .A2(_06693_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _07405_ (.A1(_06668_),
    .A2(_00425_),
    .B1(_00426_),
    .B2(_06711_),
    .C(_05171_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07406_ (.A1(_05387_),
    .A2(_00424_),
    .B(_00427_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07407_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-23] ),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07408_ (.A1(_05409_),
    .A2(_05474_),
    .B(_05518_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07409_ (.A1(_06232_),
    .A2(_06645_),
    .B(_05442_),
    .C(_06146_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07410_ (.A1(_06146_),
    .A2(_00429_),
    .B(_00430_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07411_ (.A1(_05387_),
    .A2(_00431_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07412_ (.A1(_05387_),
    .A2(_00428_),
    .B(_00432_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07413_ (.A1(_05507_),
    .A2(_06788_),
    .B(_00341_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07414_ (.A1(_05658_),
    .A2(_06705_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07415_ (.A1(_05658_),
    .A2(_00433_),
    .B1(_00434_),
    .B2(_06732_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07416_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-22] ),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07417_ (.A1(_06059_),
    .A2(_00435_),
    .B(_00436_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07418_ (.A1(_06232_),
    .A2(_06621_),
    .B(_06676_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07419_ (.A1(_06624_),
    .A2(_00343_),
    .B1(_00437_),
    .B2(_05658_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07420_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-21] ),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07421_ (.A1(_06059_),
    .A2(_00438_),
    .B(_00439_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07422_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-20] ),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07423_ (.A1(_05778_),
    .A2(_06754_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07424_ (.A1(_06630_),
    .A2(_00441_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07425_ (.A1(_05420_),
    .A2(_06092_),
    .B(_05561_),
    .C(_06232_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07426_ (.A1(_05409_),
    .A2(_05984_),
    .B(_06146_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07427_ (.A1(_06146_),
    .A2(_00442_),
    .B1(_00443_),
    .B2(_00444_),
    .C(_05280_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07428_ (.A1(_06059_),
    .A2(_00440_),
    .B(_00445_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07429_ (.A1(_05886_),
    .A2(_06754_),
    .B(_06646_),
    .C(_05658_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07430_ (.A1(_06232_),
    .A2(_06756_),
    .B(_06820_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07431_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-19] ),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07432_ (.A1(_05822_),
    .A2(_00446_),
    .A3(_00447_),
    .B(_00448_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07433_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-18] ),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07434_ (.A1(_05658_),
    .A2(_06830_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07435_ (.A1(_05409_),
    .A2(_05420_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07436_ (.A1(_05409_),
    .A2(_06092_),
    .B(_00451_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07437_ (.A1(_06698_),
    .A2(_00450_),
    .B1(_00452_),
    .B2(_05658_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07438_ (.A1(_05387_),
    .A2(_00453_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07439_ (.A1(_05387_),
    .A2(_00449_),
    .B(_00454_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07440_ (.A1(_06232_),
    .A2(_05940_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07441_ (.A1(_06146_),
    .A2(_05463_),
    .A3(_06125_),
    .B(_00455_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07442_ (.A1(_05409_),
    .A2(_05973_),
    .B1(_06622_),
    .B2(_06816_),
    .C(_00456_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07443_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-17] ),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07444_ (.A1(_06059_),
    .A2(_00457_),
    .B(_00458_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07445_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-16] ),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07446_ (.A1(_06713_),
    .A2(_05897_),
    .B1(_06070_),
    .B2(_06721_),
    .C(_05658_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07447_ (.A1(_06795_),
    .A2(_05995_),
    .B(_06826_),
    .C(_05658_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07448_ (.A1(_05182_),
    .A2(_00461_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07449_ (.A1(_05387_),
    .A2(_00459_),
    .B1(_00460_),
    .B2(_00462_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07450_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-15] ),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07451_ (.A1(_05518_),
    .A2(_05789_),
    .B1(_06070_),
    .B2(_06721_),
    .C(_05658_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07452_ (.A1(_05496_),
    .A2(_05713_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07453_ (.A1(_05658_),
    .A2(_06656_),
    .A3(_00465_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07454_ (.A1(_05182_),
    .A2(_00466_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07455_ (.A1(_05387_),
    .A2(_00463_),
    .B1(_00464_),
    .B2(_00467_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07456_ (.A1(_05409_),
    .A2(_06734_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07457_ (.A1(_05431_),
    .A2(_06705_),
    .B(_00468_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07458_ (.A1(_05658_),
    .A2(_00451_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07459_ (.A1(_05658_),
    .A2(_00469_),
    .B1(_00470_),
    .B2(_06711_),
    .C(_05182_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07460_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-14] ),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07461_ (.A1(_00471_),
    .A2(_00472_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07462_ (.A1(_05897_),
    .A2(_06666_),
    .B(_05409_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07463_ (.A1(_06778_),
    .A2(_06787_),
    .B(_05658_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07464_ (.A1(_06232_),
    .A2(_05572_),
    .A3(_05886_),
    .B(_06624_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07465_ (.A1(_05442_),
    .A2(_00475_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07466_ (.A1(_00473_),
    .A2(_00474_),
    .B1(_00476_),
    .B2(_05658_),
    .C(_05182_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07467_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-13] ),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07468_ (.A1(_00477_),
    .A2(_00478_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07469_ (.A1(_06713_),
    .A2(_06211_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07470_ (.A1(_05409_),
    .A2(_00425_),
    .B(_00479_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07471_ (.A1(_05409_),
    .A2(_05442_),
    .A3(_05875_),
    .B(_00480_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07472_ (.A1(_06799_),
    .A2(_00308_),
    .B1(_00481_),
    .B2(_05658_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07473_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-12] ),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07474_ (.A1(_06059_),
    .A2(_00482_),
    .B(_00483_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07475_ (.A1(_06651_),
    .A2(_06373_),
    .B1(_06754_),
    .B2(_06756_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07476_ (.A1(_05658_),
    .A2(_00484_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07477_ (.A1(_05409_),
    .A2(_05995_),
    .B1(_06221_),
    .B2(_06787_),
    .C(_06146_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07478_ (.A1(_05171_),
    .A2(_00485_),
    .A3(_00486_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07479_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-11] ),
    .B(_00487_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07480_ (.I(_00488_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07481_ (.A1(_05583_),
    .A2(_06754_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07482_ (.A1(_00450_),
    .A2(_00489_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07483_ (.A1(_05658_),
    .A2(_05529_),
    .A3(_06651_),
    .A4(_06712_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07484_ (.A1(_05182_),
    .A2(_00490_),
    .A3(_00491_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07485_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-10] ),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07486_ (.A1(_00492_),
    .A2(_00493_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07487_ (.A1(_05995_),
    .A2(_06221_),
    .B(_06146_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07488_ (.A1(_06753_),
    .A2(_06789_),
    .B(_00494_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07489_ (.A1(_06232_),
    .A2(_06070_),
    .B(_00455_),
    .C(_05658_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07490_ (.A1(_06703_),
    .A2(_00496_),
    .B(_05182_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07491_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07492_ (.A1(_00495_),
    .A2(_00497_),
    .B(_00498_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07493_ (.A1(_06790_),
    .A2(_06827_),
    .B1(_00455_),
    .B2(_06797_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07494_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-8] ),
    .I1(_00499_),
    .S(_00395_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07495_ (.I(_00500_),
    .Z(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07496_ (.A1(_06232_),
    .A2(_06713_),
    .A3(_05897_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07497_ (.A1(_06146_),
    .A2(_05745_),
    .A3(_00501_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07498_ (.A1(_05658_),
    .A2(_05724_),
    .A3(_06761_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07499_ (.A1(_05171_),
    .A2(_00503_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07500_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-7] ),
    .B1(_00502_),
    .B2(_00504_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07501_ (.I(_00505_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07502_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-6] ),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07503_ (.A1(_05409_),
    .A2(_05995_),
    .B(_06761_),
    .C(_06146_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07504_ (.A1(_05431_),
    .A2(_06779_),
    .B(_00455_),
    .C(_05658_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07505_ (.A1(_05182_),
    .A2(_00507_),
    .A3(_00508_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07506_ (.A1(_05387_),
    .A2(_00506_),
    .B(_00509_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07507_ (.A1(_06726_),
    .A2(_06806_),
    .B(_05658_),
    .C(_05474_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07508_ (.A1(_06146_),
    .A2(_05897_),
    .B(_05182_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07509_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07510_ (.A1(_00510_),
    .A2(_00511_),
    .B(_00512_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07511_ (.A1(_06703_),
    .A2(_06629_),
    .B(_06766_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07512_ (.A1(_05409_),
    .A2(_06458_),
    .B1(_00347_),
    .B2(_06753_),
    .C(_05658_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07513_ (.A1(_05658_),
    .A2(_00513_),
    .B(_00514_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07514_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-4] ),
    .I1(_00515_),
    .S(_00395_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07515_ (.I(_00516_),
    .Z(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07516_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-3] ),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07517_ (.A1(_05875_),
    .A2(_06666_),
    .B(_06613_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07518_ (.A1(_05713_),
    .A2(_06614_),
    .B(_00518_),
    .C(_05658_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07519_ (.A1(_05658_),
    .A2(_06623_),
    .A3(_00465_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07520_ (.A1(_05182_),
    .A2(_00520_),
    .ZN(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07521_ (.A1(_05387_),
    .A2(_00517_),
    .B1(_00519_),
    .B2(_00521_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07522_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-2] ),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07523_ (.A1(_05940_),
    .A2(_06622_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07524_ (.A1(_00419_),
    .A2(_00523_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07525_ (.A1(_05658_),
    .A2(_06651_),
    .A3(_06733_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _07526_ (.A1(_05658_),
    .A2(_00524_),
    .B1(_00525_),
    .B2(_00330_),
    .C(_05171_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07527_ (.A1(_05387_),
    .A2(_00522_),
    .B(_00526_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07528_ (.A1(_05409_),
    .A2(_06715_),
    .B(_06566_),
    .C(_06146_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07529_ (.A1(_05496_),
    .A2(_06806_),
    .B(_05908_),
    .C(_05658_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07530_ (.A1(_05171_),
    .A2(_00527_),
    .A3(_00528_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07531_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-1] ),
    .B(_00529_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07532_ (.I(_00530_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07533_ (.A1(_05409_),
    .A2(_05420_),
    .A3(_06092_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07534_ (.A1(_06232_),
    .A2(_05897_),
    .B(_05658_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07535_ (.A1(_06645_),
    .A2(_06748_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07536_ (.A1(_06232_),
    .A2(_05919_),
    .B(_00533_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07537_ (.A1(_00531_),
    .A2(_00532_),
    .B1(_00534_),
    .B2(_05658_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07538_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ),
    .I1(_00535_),
    .S(_00395_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07539_ (.I(_00536_),
    .Z(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07540_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[1] ),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07541_ (.A1(_05778_),
    .A2(_06721_),
    .B(_06373_),
    .C(_05658_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07542_ (.A1(_05658_),
    .A2(_05529_),
    .A3(_00441_),
    .A4(_00443_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07543_ (.A1(_05182_),
    .A2(_00539_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07544_ (.A1(_05387_),
    .A2(_00537_),
    .B1(_00538_),
    .B2(_00540_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07545_ (.A1(_05572_),
    .A2(_05550_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07546_ (.A1(_05409_),
    .A2(_00541_),
    .B(_06682_),
    .C(_06146_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07547_ (.A1(_05951_),
    .A2(_06704_),
    .B(_00479_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07548_ (.A1(_05658_),
    .A2(_06661_),
    .A3(_00543_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07549_ (.A1(_05182_),
    .A2(_00542_),
    .A3(_00544_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07550_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[2] ),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07551_ (.A1(_00545_),
    .A2(_00546_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07552_ (.A1(_05550_),
    .A2(_06789_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07553_ (.A1(_06092_),
    .A2(_06622_),
    .B(_00547_),
    .C(_05658_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07554_ (.A1(_00348_),
    .A2(_06733_),
    .A3(_06756_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07555_ (.A1(_05182_),
    .A2(_00548_),
    .A3(_00549_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07556_ (.A1(_05822_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[3] ),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07557_ (.A1(_00550_),
    .A2(_00551_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07558_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[4] ),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07559_ (.I(_00350_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07560_ (.A1(_05409_),
    .A2(_05594_),
    .B(_06735_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07561_ (.A1(_06059_),
    .A2(_00552_),
    .B1(_00553_),
    .B2(_00554_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07562_ (.A1(_05409_),
    .A2(_00541_),
    .B(_06693_),
    .C(_05658_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07563_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[5] ),
    .I1(_00555_),
    .S(_00395_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07564_ (.I(_00556_),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07565_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[16] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-15] ),
    .S(_00395_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07566_ (.I(_00557_),
    .Z(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07567_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[17] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-14] ),
    .S(_00395_),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07568_ (.I(_00558_),
    .Z(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07569_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[18] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ),
    .S(_00395_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07570_ (.I(_00559_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07571_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[19] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-12] ),
    .S(_00395_),
    .Z(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07572_ (.I(_00560_),
    .Z(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07573_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[20] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-11] ),
    .S(_00395_),
    .Z(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07574_ (.I(_00561_),
    .Z(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07575_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[21] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-10] ),
    .S(_00395_),
    .Z(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07576_ (.I(_00562_),
    .Z(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07577_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[22] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-9] ),
    .S(_00395_),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07578_ (.I(_00563_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07579_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[23] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-8] ),
    .S(_00395_),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07580_ (.I(_00564_),
    .Z(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07581_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[24] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-7] ),
    .S(_00395_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07582_ (.I(_00565_),
    .Z(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07583_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[25] ),
    .I1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-6] ),
    .S(_00395_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07584_ (.I(_00566_),
    .Z(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07585_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[26] ),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07586_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-5] ),
    .A2(_05182_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07587_ (.A1(_05387_),
    .A2(_00567_),
    .B(_00568_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07588_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[27] ),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07589_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-4] ),
    .A2(_05182_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07590_ (.A1(_05387_),
    .A2(_00569_),
    .B(_00570_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07591_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[28] ),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07592_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-3] ),
    .A2(_05182_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07593_ (.A1(_05387_),
    .A2(_00571_),
    .B(_00572_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07594_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[29] ),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07595_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-2] ),
    .A2(_05182_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07596_ (.A1(_05387_),
    .A2(_00573_),
    .B(_00574_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07597_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[30] ),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07598_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-1] ),
    .A2(_05182_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07599_ (.A1(_05387_),
    .A2(_00575_),
    .B(_00576_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07600_ (.I(\DDS_Stage.LCU.SelMuxConfigReg ),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07601_ (.I(_00577_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07602_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-15] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-15] ),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07603_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-15] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-15] ),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07604_ (.A1(_00578_),
    .A2(_00580_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07605_ (.A1(\DDS_Stage.xPoints_Generator1.CosNew[-15] ),
    .A2(_00578_),
    .B1(_00579_),
    .B2(_00581_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07606_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-15] ),
    .A2(_05280_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07607_ (.A1(_06059_),
    .A2(_00582_),
    .B(_00583_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07608_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-14] ),
    .A2(_05822_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07609_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-14] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-14] ),
    .A3(_00579_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07610_ (.A1(_00577_),
    .A2(_00585_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07611_ (.A1(_00577_),
    .A2(\DDS_Stage.xPoints_Generator1.CosNew[-14] ),
    .B(_05182_),
    .C(_00586_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07612_ (.A1(_00584_),
    .A2(_00587_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07613_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-14] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-14] ),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07614_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-14] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-14] ),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07615_ (.A1(_00579_),
    .A2(_00588_),
    .B(_00589_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07616_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-13] ),
    .A3(_00590_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07617_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-13] ),
    .I1(_00591_),
    .S(_00577_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07618_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ),
    .I1(_00592_),
    .S(_00395_),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07619_ (.I(_00593_),
    .Z(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07620_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-13] ),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07621_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-13] ),
    .B(_00590_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07622_ (.A1(_00594_),
    .A2(_00595_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07623_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-12] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-12] ),
    .A3(_00596_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07624_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-12] ),
    .I1(_00597_),
    .S(_00577_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07625_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-12] ),
    .I1(_00598_),
    .S(_00395_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07626_ (.I(_00599_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07627_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-12] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-12] ),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07628_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-12] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-12] ),
    .B(_00596_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07629_ (.A1(_00600_),
    .A2(_00601_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07630_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-11] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-11] ),
    .A3(_00602_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07631_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-11] ),
    .I1(_00603_),
    .S(_00577_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07632_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-11] ),
    .I1(_00604_),
    .S(_00395_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07633_ (.I(_00605_),
    .Z(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07634_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-11] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-11] ),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07635_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-11] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-11] ),
    .B(_00602_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07636_ (.A1(_00606_),
    .A2(_00607_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07637_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-10] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-10] ),
    .A3(_00608_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07638_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-10] ),
    .I1(_00609_),
    .S(_00577_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07639_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-10] ),
    .I1(_00610_),
    .S(_00395_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07640_ (.I(_00611_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07641_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-10] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-10] ),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07642_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-10] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-10] ),
    .B(_00608_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07643_ (.A1(_00612_),
    .A2(_00613_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07644_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-9] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-9] ),
    .A3(_00614_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07645_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-9] ),
    .I1(_00615_),
    .S(_00577_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07646_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-9] ),
    .I1(_00616_),
    .S(_00395_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07647_ (.I(_00617_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07648_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-9] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-9] ),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07649_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-9] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-9] ),
    .B(_00614_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07650_ (.A1(_00618_),
    .A2(_00619_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07651_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-8] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-8] ),
    .A3(_00620_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07652_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-8] ),
    .I1(_00621_),
    .S(_00577_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07653_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-8] ),
    .I1(_00622_),
    .S(_00395_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07654_ (.I(_00623_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07655_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-8] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-8] ),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07656_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-8] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-8] ),
    .B(_00620_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07657_ (.A1(_00624_),
    .A2(_00625_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07658_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-7] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-7] ),
    .A3(_00626_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07659_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-7] ),
    .I1(_00627_),
    .S(_00577_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07660_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-7] ),
    .I1(_00628_),
    .S(_00395_),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07661_ (.I(_00629_),
    .Z(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07662_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-7] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-7] ),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07663_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-7] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-7] ),
    .B(_00626_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07664_ (.A1(_00630_),
    .A2(_00631_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07665_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-6] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-6] ),
    .A3(_00632_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07666_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-6] ),
    .I1(_00633_),
    .S(_00577_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07667_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-6] ),
    .I1(_00634_),
    .S(_00395_),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07668_ (.I(_00635_),
    .Z(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07669_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-6] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-6] ),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07670_ (.A1(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-6] ),
    .A2(\DDS_Stage.xPoints_Generator1.RegFrequency[-6] ),
    .B(_00632_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07671_ (.A1(_00636_),
    .A2(_00637_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07672_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-5] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-5] ),
    .A3(_00638_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07673_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-5] ),
    .I1(_00639_),
    .S(_00577_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07674_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-5] ),
    .I1(_00640_),
    .S(_00395_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07675_ (.I(_00641_),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07676_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-5] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-5] ),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07677_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-5] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-5] ),
    .B(_00638_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07678_ (.A1(_00642_),
    .A2(_00643_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07679_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-4] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-4] ),
    .A3(_00644_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07680_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-4] ),
    .I1(_00645_),
    .S(_00577_),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07681_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-4] ),
    .I1(_00646_),
    .S(_00395_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07682_ (.I(_00647_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07683_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-4] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-4] ),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07684_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-4] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-4] ),
    .B(_00644_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07685_ (.A1(_00648_),
    .A2(_00649_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07686_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-3] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-3] ),
    .A3(_00650_),
    .Z(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07687_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-3] ),
    .I1(_00651_),
    .S(_00577_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07688_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-3] ),
    .I1(_00652_),
    .S(_00395_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07689_ (.I(_00653_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07690_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-3] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-3] ),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07691_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-3] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-3] ),
    .B(_00650_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07692_ (.A1(_00654_),
    .A2(_00655_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07693_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-2] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-2] ),
    .A3(_00656_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07694_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-2] ),
    .I1(_00657_),
    .S(_00577_),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07695_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-2] ),
    .I1(_00658_),
    .S(_00395_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07696_ (.I(_00659_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07697_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-2] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-2] ),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07698_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-2] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-2] ),
    .B(_00656_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07699_ (.A1(_00660_),
    .A2(_00661_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07700_ (.A1(\DDS_Stage.xPoints_Generator1.RegFrequency[-1] ),
    .A2(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-1] ),
    .A3(_00662_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07701_ (.I0(\DDS_Stage.xPoints_Generator1.CosNew[-1] ),
    .I1(_00663_),
    .S(_00577_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07702_ (.I0(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-1] ),
    .I1(_00664_),
    .S(_00395_),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07703_ (.I(_00665_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07704_ (.A1(net36),
    .A2(_05237_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07705_ (.I(_00666_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07706_ (.I0(net2),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-15] ),
    .S(_00667_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07707_ (.I(_00668_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07708_ (.I0(net8),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-14] ),
    .S(_00667_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07709_ (.I(_00669_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07710_ (.I0(net114),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-13] ),
    .S(_00667_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07711_ (.I(_00670_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07712_ (.I0(net10),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-12] ),
    .S(_00667_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07713_ (.I(_00671_),
    .Z(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07714_ (.I0(net118),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-11] ),
    .S(_00667_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07715_ (.I(_00672_),
    .Z(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07716_ (.I0(net112),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-10] ),
    .S(_00667_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07717_ (.I(_00673_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07718_ (.I0(net116),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-9] ),
    .S(_00667_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07719_ (.I(_00674_),
    .Z(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07720_ (.I0(net104),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-8] ),
    .S(_00667_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07721_ (.I(_00675_),
    .Z(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07722_ (.I0(net108),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-7] ),
    .S(_00667_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07723_ (.I(_00676_),
    .Z(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07724_ (.I0(net106),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-6] ),
    .S(_00667_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07725_ (.I(_00677_),
    .Z(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07726_ (.I0(net110),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-5] ),
    .S(_00667_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07727_ (.I(_00678_),
    .Z(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07728_ (.I0(net4),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-4] ),
    .S(_00667_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07729_ (.I(_00679_),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07730_ (.I0(net5),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-3] ),
    .S(_00667_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07731_ (.I(_00680_),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07732_ (.I0(net6),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-2] ),
    .S(_00667_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07733_ (.I(_00681_),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07734_ (.I0(net7),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-1] ),
    .S(_00667_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07735_ (.I(_00682_),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07736_ (.A1(net36),
    .A2(_05324_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07737_ (.I(_00683_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07738_ (.I0(net2),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-15] ),
    .S(_00684_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07739_ (.I(_00685_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07740_ (.I0(net8),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-14] ),
    .S(_00684_),
    .Z(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07741_ (.I(_00686_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07742_ (.I0(net114),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-13] ),
    .S(_00684_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07743_ (.I(_00687_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07744_ (.I0(net120),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-12] ),
    .S(_00684_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07745_ (.I(_00688_),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07746_ (.I0(net118),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-11] ),
    .S(_00684_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07747_ (.I(_00689_),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07748_ (.I0(net112),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-10] ),
    .S(_00684_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07749_ (.I(_00690_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07750_ (.I0(net116),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-9] ),
    .S(_00684_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07751_ (.I(_00691_),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07752_ (.I0(net104),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-8] ),
    .S(_00684_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07753_ (.I(_00692_),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07754_ (.I0(net108),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-7] ),
    .S(_00684_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07755_ (.I(_00693_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07756_ (.I0(net106),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-6] ),
    .S(_00684_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07757_ (.I(_00694_),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07758_ (.I0(net110),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-5] ),
    .S(_00684_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07759_ (.I(_00695_),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07760_ (.I0(net4),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-4] ),
    .S(_00684_),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07761_ (.I(_00696_),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07762_ (.I0(net5),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-3] ),
    .S(_00684_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07763_ (.I(_00697_),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07764_ (.I0(net6),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-2] ),
    .S(_00684_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07765_ (.I(_00698_),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07766_ (.I0(net7),
    .I1(\DDS_Stage.xPoints_Generator1.RegP[-1] ),
    .S(_00684_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07767_ (.I(_00699_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07768_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-15] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-15] ),
    .S(_00402_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07769_ (.I(_00700_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07770_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-14] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-14] ),
    .S(_00402_),
    .Z(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07771_ (.I(_00701_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07772_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-13] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-13] ),
    .S(_00402_),
    .Z(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07773_ (.I(_00702_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07774_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-12] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-12] ),
    .S(_00402_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07775_ (.I(_00703_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07776_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-11] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-11] ),
    .S(_00402_),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07777_ (.I(_00704_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07778_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-10] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-10] ),
    .S(_00402_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07779_ (.I(_00705_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07780_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-9] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-9] ),
    .S(_00402_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07781_ (.I(_00706_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07782_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-8] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-8] ),
    .S(_00402_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07783_ (.I(_00707_),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07784_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-7] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-7] ),
    .S(_00402_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07785_ (.I(_00708_),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07786_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-6] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-6] ),
    .S(_00402_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07787_ (.I(_00709_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07788_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-5] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-5] ),
    .S(_00402_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07789_ (.I(_00710_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07790_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-4] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-4] ),
    .S(_00402_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07791_ (.I(_00711_),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07792_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-3] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-3] ),
    .S(_00402_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07793_ (.I(_00712_),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07794_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-2] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-2] ),
    .S(_00402_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07795_ (.I(_00713_),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07796_ (.I0(\DDS_Stage.xPoints_Generator1.RegFrequency[-1] ),
    .I1(\DDS_Stage.xPoints_Generator1.RegF[-1] ),
    .S(_00402_),
    .Z(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07797_ (.I(_00714_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07798_ (.I0(net58),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[16] ),
    .S(_00395_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07799_ (.I(_00715_),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07800_ (.I0(_00355_),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[17] ),
    .S(_00395_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07801_ (.I(_00716_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07802_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[18] ),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07803_ (.A1(_05387_),
    .A2(_00358_),
    .B(_00717_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07804_ (.I0(net60),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[19] ),
    .S(_00395_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07805_ (.I(_00718_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07806_ (.I0(net61),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[20] ),
    .S(_00395_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07807_ (.I(_00719_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07808_ (.I0(_00370_),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[21] ),
    .S(_00395_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07809_ (.I(_00720_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07810_ (.I0(_00373_),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[22] ),
    .S(_00395_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07811_ (.I(_00721_),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07812_ (.I0(_00376_),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[23] ),
    .S(_00395_),
    .Z(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07813_ (.I(_00722_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07814_ (.I0(_00379_),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[24] ),
    .S(_00395_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07815_ (.I(_00723_),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07816_ (.I0(_00382_),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[25] ),
    .S(_00395_),
    .Z(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07817_ (.I(_00724_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07818_ (.A1(_05280_),
    .A2(_00385_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07819_ (.A1(_06059_),
    .A2(_00567_),
    .B(_00725_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07820_ (.A1(_05280_),
    .A2(_00388_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07821_ (.A1(_06059_),
    .A2(_00569_),
    .B(_00726_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07822_ (.A1(_05280_),
    .A2(net63),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07823_ (.A1(_06059_),
    .A2(_00571_),
    .B(_00727_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07824_ (.A1(_05280_),
    .A2(_00394_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07825_ (.A1(_06059_),
    .A2(_00573_),
    .B(_00728_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07826_ (.A1(_05280_),
    .A2(_00398_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07827_ (.A1(_06059_),
    .A2(_00575_),
    .B(_00729_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07828_ (.A1(net155),
    .A2(_00373_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07829_ (.A1(_06308_),
    .A2(_00379_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07830_ (.A1(net152),
    .A2(_00376_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07831_ (.A1(_00731_),
    .A2(_00732_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07832_ (.A1(_00731_),
    .A2(_00732_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07833_ (.A1(_00733_),
    .A2(_00734_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07834_ (.A1(_00730_),
    .A2(_00735_),
    .B(_00733_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07835_ (.A1(_00730_),
    .A2(_00735_),
    .Z(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07836_ (.A1(_05833_),
    .A2(_05398_),
    .A3(_00388_),
    .A4(_00385_),
    .Z(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07837_ (.A1(_05864_),
    .A2(_00382_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07838_ (.A1(_05398_),
    .A2(_00388_),
    .B1(_00385_),
    .B2(_05833_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07839_ (.A1(_00738_),
    .A2(_00739_),
    .A3(_00740_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07840_ (.A1(_00738_),
    .A2(_00741_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07841_ (.A1(_06179_),
    .A2(_00382_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07842_ (.A1(_05864_),
    .A2(_05833_),
    .A3(_00388_),
    .A4(_00385_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07843_ (.A1(_05833_),
    .A2(_00388_),
    .B1(_00385_),
    .B2(_05864_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07844_ (.A1(_00744_),
    .A2(_00745_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07845_ (.A1(_00743_),
    .A2(_00746_),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07846_ (.A1(_00742_),
    .A2(_00747_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07847_ (.A1(_00737_),
    .A2(_00748_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07848_ (.A1(net152),
    .A2(_00373_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07849_ (.A1(_06308_),
    .A2(_00376_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07850_ (.A1(_06179_),
    .A2(_00379_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07851_ (.A1(_00751_),
    .A2(_00752_),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07852_ (.A1(_00751_),
    .A2(_00752_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07853_ (.A1(_00753_),
    .A2(_00754_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07854_ (.A1(_00750_),
    .A2(_00755_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07855_ (.A1(_05833_),
    .A2(_05398_),
    .A3(_00385_),
    .A4(_00382_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07856_ (.A1(_00738_),
    .A2(_00740_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07857_ (.A1(_00739_),
    .A2(_00758_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07858_ (.A1(_00757_),
    .A2(_00759_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07859_ (.A1(_00757_),
    .A2(_00759_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07860_ (.A1(_00756_),
    .A2(_00760_),
    .B(_00761_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07861_ (.A1(_00749_),
    .A2(_00762_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07862_ (.A1(_00736_),
    .A2(_00763_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07863_ (.A1(_06618_),
    .A2(_00370_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07864_ (.A1(_00764_),
    .A2(_00765_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07865_ (.A1(_00736_),
    .A2(_00763_),
    .B(_00766_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07866_ (.I(_00767_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07867_ (.A1(_00764_),
    .A2(_00765_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07868_ (.A1(_00749_),
    .A2(_00762_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07869_ (.A1(net137),
    .A2(_00355_),
    .A3(_06633_),
    .A4(_06627_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07870_ (.A1(net58),
    .A2(_06633_),
    .B1(_06627_),
    .B2(_00355_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07871_ (.I(_00772_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07872_ (.A1(_00773_),
    .A2(_00771_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07873_ (.A1(_00357_),
    .A2(_06598_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07874_ (.A1(net92),
    .A2(net153),
    .B1(_06523_),
    .B2(net143),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07875_ (.A1(net92),
    .A2(net143),
    .A3(_06416_),
    .A4(net156),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07876_ (.A1(_00775_),
    .A2(_00776_),
    .B(_00777_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07877_ (.A1(_00357_),
    .A2(_06618_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07878_ (.A1(_00367_),
    .A2(_06523_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07879_ (.A1(_00363_),
    .A2(_06598_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07880_ (.A1(_00779_),
    .A2(_00780_),
    .A3(_00781_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07881_ (.A1(_00782_),
    .A2(_00778_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07882_ (.A1(net157),
    .A2(_00782_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07883_ (.A1(_00774_),
    .A2(_00783_),
    .B(_00784_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07884_ (.A1(_06637_),
    .A2(net58),
    .B1(_00355_),
    .B2(_06633_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07885_ (.I(_00786_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07886_ (.A1(_06637_),
    .A2(net58),
    .A3(_00355_),
    .A4(_06633_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07887_ (.A1(_00787_),
    .A2(_00788_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07888_ (.A1(net91),
    .A2(net156),
    .B1(_06598_),
    .B2(net142),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07889_ (.A1(net91),
    .A2(net142),
    .A3(net156),
    .A4(_06598_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07890_ (.A1(_00779_),
    .A2(_00790_),
    .B(_00791_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07891_ (.A1(_00357_),
    .A2(_06627_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07892_ (.A1(net158),
    .A2(_06598_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07893_ (.A1(net143),
    .A2(_06618_),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07894_ (.A1(_00793_),
    .A2(_00794_),
    .A3(_00795_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07895_ (.A1(_00792_),
    .A2(_00796_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07896_ (.A1(_00789_),
    .A2(_00797_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07897_ (.A1(_00785_),
    .A2(_00798_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07898_ (.A1(_00785_),
    .A2(_00798_),
    .ZN(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07899_ (.A1(_00771_),
    .A2(_00799_),
    .B(_00800_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07900_ (.A1(_00792_),
    .A2(_00796_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07901_ (.A1(_00789_),
    .A2(_00797_),
    .B(_00802_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07902_ (.A1(net91),
    .A2(_06598_),
    .B1(_06618_),
    .B2(net143),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07903_ (.A1(net91),
    .A2(net142),
    .A3(_06598_),
    .A4(_06618_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07904_ (.A1(_00793_),
    .A2(_00804_),
    .B(_00805_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07905_ (.A1(_00357_),
    .A2(_06633_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07906_ (.A1(_00367_),
    .A2(_06618_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07907_ (.A1(_00363_),
    .A2(_06627_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07908_ (.A1(_00807_),
    .A2(_00808_),
    .A3(_00809_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07909_ (.A1(_00806_),
    .A2(_00810_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07910_ (.A1(_06637_),
    .A2(_00355_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07911_ (.A1(_06642_),
    .A2(_00352_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07912_ (.A1(_00391_),
    .A2(_05398_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07913_ (.A1(_00813_),
    .A2(_00814_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07914_ (.A1(_00812_),
    .A2(_00815_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07915_ (.A1(_00811_),
    .A2(_00816_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07916_ (.A1(_00803_),
    .A2(_00817_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07917_ (.A1(_00788_),
    .A2(_00818_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07918_ (.A1(_00801_),
    .A2(_00819_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07919_ (.A1(_00801_),
    .A2(_00819_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07920_ (.A1(_00770_),
    .A2(_00820_),
    .B(_00821_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07921_ (.A1(_06598_),
    .A2(_00373_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07922_ (.A1(net152),
    .A2(_00379_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07923_ (.A1(net155),
    .A2(_00376_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07924_ (.A1(_00824_),
    .A2(_00825_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07925_ (.A1(_00823_),
    .A2(_00826_),
    .Z(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07926_ (.A1(_05864_),
    .A2(_05833_),
    .A3(_00388_),
    .A4(_00385_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07927_ (.A1(_00743_),
    .A2(_00745_),
    .B(_00828_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07928_ (.I(_00829_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07929_ (.A1(_06308_),
    .A2(_00382_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07930_ (.A1(_06179_),
    .A2(_05864_),
    .A3(_00388_),
    .A4(_00385_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07931_ (.A1(_05864_),
    .A2(_00388_),
    .B1(_00385_),
    .B2(_06179_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07932_ (.A1(_00832_),
    .A2(_00833_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07933_ (.A1(_00831_),
    .A2(_00834_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07934_ (.A1(_00830_),
    .A2(_00835_),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07935_ (.A1(_00827_),
    .A2(_00836_),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07936_ (.A1(_00737_),
    .A2(_00748_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07937_ (.A1(_00742_),
    .A2(_00747_),
    .B(_00838_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07938_ (.A1(_00837_),
    .A2(_00839_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07939_ (.A1(_00803_),
    .A2(_00817_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07940_ (.A1(_00788_),
    .A2(_00818_),
    .B(_00841_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07941_ (.A1(_06637_),
    .A2(_00355_),
    .A3(_00815_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07942_ (.A1(_00813_),
    .A2(_00814_),
    .B(_00843_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07943_ (.A1(_00394_),
    .A2(_05398_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07944_ (.A1(_00844_),
    .A2(_00845_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07945_ (.A1(_00806_),
    .A2(_00810_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07946_ (.A1(_00811_),
    .A2(_00816_),
    .B(_00847_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07947_ (.A1(net142),
    .A2(_06627_),
    .B1(_06618_),
    .B2(net92),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07948_ (.A1(net92),
    .A2(net142),
    .A3(_06627_),
    .A4(_06618_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07949_ (.A1(_00807_),
    .A2(_00849_),
    .B(_00850_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07950_ (.A1(_00357_),
    .A2(_06637_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07951_ (.A1(net74),
    .A2(_06627_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07952_ (.A1(net143),
    .A2(_06633_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07953_ (.A1(_00852_),
    .A2(_00853_),
    .A3(_00854_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07954_ (.A1(_00851_),
    .A2(_00855_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07955_ (.A1(_06642_),
    .A2(_00355_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07956_ (.A1(_06649_),
    .A2(_00352_),
    .A3(_00391_),
    .A4(_05833_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07957_ (.A1(_06649_),
    .A2(net138),
    .B1(_00391_),
    .B2(_05833_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07958_ (.A1(_00858_),
    .A2(_00859_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07959_ (.A1(_00857_),
    .A2(_00860_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07960_ (.A1(_00856_),
    .A2(_00861_),
    .Z(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07961_ (.A1(_00848_),
    .A2(_00862_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07962_ (.A1(_00846_),
    .A2(_00863_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07963_ (.A1(_00842_),
    .A2(_00864_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07964_ (.A1(_00840_),
    .A2(_00865_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07965_ (.A1(_00822_),
    .A2(_00866_),
    .Z(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07966_ (.A1(_00822_),
    .A2(_00866_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07967_ (.A1(_00769_),
    .A2(_00867_),
    .B(_00868_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07968_ (.A1(_00837_),
    .A2(_00839_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07969_ (.A1(_00824_),
    .A2(_00825_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07970_ (.A1(_00823_),
    .A2(_00826_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07971_ (.A1(_00871_),
    .A2(_00872_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07972_ (.A1(_00870_),
    .A2(_00873_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07973_ (.A1(_06627_),
    .A2(_00370_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07974_ (.A1(_00874_),
    .A2(_00875_),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07975_ (.A1(_00842_),
    .A2(_00864_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07976_ (.A1(_00840_),
    .A2(_00865_),
    .B(_00877_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07977_ (.A1(_00848_),
    .A2(_00862_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07978_ (.A1(_00846_),
    .A2(_00863_),
    .B(_00879_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07979_ (.A1(_00857_),
    .A2(_00860_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07980_ (.A1(_00858_),
    .A2(_00881_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07981_ (.A1(_00394_),
    .A2(_05833_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07982_ (.A1(_00398_),
    .A2(_05398_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07983_ (.A1(_00883_),
    .A2(_00884_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07984_ (.A1(_00883_),
    .A2(_00884_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07985_ (.A1(_00885_),
    .A2(_00886_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07986_ (.A1(_00882_),
    .A2(_00887_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07987_ (.A1(_00851_),
    .A2(_00855_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07988_ (.A1(_00856_),
    .A2(_00861_),
    .B(_00889_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07989_ (.A1(_00363_),
    .A2(_06633_),
    .B1(_06627_),
    .B2(net91),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07990_ (.A1(net91),
    .A2(_00363_),
    .A3(_06633_),
    .A4(_06627_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07991_ (.A1(_00852_),
    .A2(_00891_),
    .B(_00892_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07992_ (.A1(_06642_),
    .A2(_00357_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07993_ (.A1(net74),
    .A2(_06633_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07994_ (.A1(_00363_),
    .A2(_06637_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07995_ (.A1(_00894_),
    .A2(_00895_),
    .A3(_00896_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07996_ (.A1(_00897_),
    .A2(_00893_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07997_ (.A1(_06649_),
    .A2(_00355_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _07998_ (.A1(_06654_),
    .A2(_00352_),
    .A3(_00391_),
    .A4(_05864_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07999_ (.A1(_06654_),
    .A2(_00352_),
    .B1(_00391_),
    .B2(_05864_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08000_ (.A1(_00900_),
    .A2(_00901_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08001_ (.A1(_00899_),
    .A2(_00902_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08002_ (.A1(_00903_),
    .A2(_00898_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08003_ (.A1(_00904_),
    .A2(_00890_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08004_ (.A1(_00888_),
    .A2(_00905_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08005_ (.A1(_00880_),
    .A2(_00906_),
    .Z(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08006_ (.A1(_00827_),
    .A2(_00836_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08007_ (.A1(_00830_),
    .A2(_00835_),
    .B(_00908_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08008_ (.A1(_00394_),
    .A2(_05398_),
    .A3(_00844_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08009_ (.A1(_00831_),
    .A2(_00832_),
    .A3(_00833_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08010_ (.A1(_00832_),
    .A2(_00911_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08011_ (.A1(_06416_),
    .A2(_00382_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08012_ (.A1(_06179_),
    .A2(_00388_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08013_ (.A1(_06308_),
    .A2(_00385_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08014_ (.A1(_00913_),
    .A2(_00914_),
    .A3(_00915_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08015_ (.A1(_00912_),
    .A2(_00916_),
    .Z(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08016_ (.A1(_06618_),
    .A2(_00373_),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08017_ (.A1(net156),
    .A2(_00379_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08018_ (.A1(_06598_),
    .A2(_00376_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08019_ (.A1(_00919_),
    .A2(_00920_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08020_ (.A1(_00918_),
    .A2(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08021_ (.A1(_00917_),
    .A2(_00922_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08022_ (.A1(_00910_),
    .A2(_00923_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08023_ (.A1(_00909_),
    .A2(_00924_),
    .Z(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08024_ (.A1(_00907_),
    .A2(_00925_),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08025_ (.A1(_00878_),
    .A2(_00926_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08026_ (.A1(_00927_),
    .A2(_00876_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08027_ (.A1(_00928_),
    .A2(_00869_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08028_ (.A1(_00929_),
    .A2(_00768_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08029_ (.A1(_05398_),
    .A2(_00385_),
    .B1(_00382_),
    .B2(_05833_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08030_ (.I(_00931_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08031_ (.A1(_00757_),
    .A2(_00932_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08032_ (.A1(_06308_),
    .A2(_00373_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08033_ (.A1(_06179_),
    .A2(_00376_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08034_ (.A1(_05864_),
    .A2(_00379_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08035_ (.A1(_00934_),
    .A2(_00935_),
    .A3(_00936_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08036_ (.A1(_00933_),
    .A2(_00937_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08037_ (.A1(_00757_),
    .A2(_00759_),
    .A3(_00756_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08038_ (.A1(_00938_),
    .A2(_00939_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08039_ (.A1(_00750_),
    .A2(_00755_),
    .B(_00753_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08040_ (.A1(_00940_),
    .A2(_00941_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08041_ (.A1(_06598_),
    .A2(_00370_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08042_ (.A1(_00938_),
    .A2(_00939_),
    .A3(_00941_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08043_ (.A1(_00942_),
    .A2(_00943_),
    .B(_00944_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08044_ (.A1(_00942_),
    .A2(_00943_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08045_ (.I(_00946_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08046_ (.A1(_00938_),
    .A2(_00939_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08047_ (.A1(net138),
    .A2(_06627_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08048_ (.A1(_00355_),
    .A2(_06618_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08049_ (.A1(_00949_),
    .A2(_00950_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08050_ (.A1(_00949_),
    .A2(_00950_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08051_ (.A1(_00952_),
    .A2(_00951_),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08052_ (.A1(net73),
    .A2(_06523_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08053_ (.A1(net92),
    .A2(_06308_),
    .B1(_06416_),
    .B2(_00363_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08054_ (.A1(net92),
    .A2(net143),
    .A3(_06308_),
    .A4(net153),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08055_ (.A1(_00954_),
    .A2(_00955_),
    .B(_00956_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08056_ (.A1(_00367_),
    .A2(_06416_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08057_ (.A1(_06523_),
    .A2(_00362_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08058_ (.A1(_00958_),
    .A2(_00959_),
    .A3(_00775_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08059_ (.A1(_00957_),
    .A2(_00960_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08060_ (.A1(_00957_),
    .A2(net85),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08061_ (.A1(_00953_),
    .A2(_00961_),
    .B(_00962_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08062_ (.A1(_00774_),
    .A2(_00783_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08063_ (.A1(_00964_),
    .A2(_00963_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08064_ (.A1(_00963_),
    .A2(net72),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08065_ (.A1(_00951_),
    .A2(_00965_),
    .B(_00966_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08066_ (.A1(_00771_),
    .A2(_00799_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08067_ (.A1(_00967_),
    .A2(_00968_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08068_ (.A1(_00967_),
    .A2(_00968_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08069_ (.A1(_00948_),
    .A2(_00969_),
    .B(_00970_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08070_ (.A1(_00770_),
    .A2(_00820_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08071_ (.A1(_00971_),
    .A2(_00972_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08072_ (.A1(_00948_),
    .A2(_00969_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08073_ (.A1(_00970_),
    .A2(_00974_),
    .B(_00972_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08074_ (.A1(_00947_),
    .A2(_00973_),
    .B(_00975_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08075_ (.A1(_00769_),
    .A2(_00867_),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08076_ (.A1(_00976_),
    .A2(_00977_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08077_ (.A1(_00976_),
    .A2(_00977_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08078_ (.A1(_00945_),
    .A2(_00978_),
    .B(_00979_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08079_ (.A1(_00930_),
    .A2(_00980_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08080_ (.A1(_05833_),
    .A2(_05398_),
    .A3(_00376_),
    .A4(_00373_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08081_ (.A1(_06179_),
    .A2(_00370_),
    .A3(_00982_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _08082_ (.A1(_06179_),
    .A2(_00370_),
    .A3(_00982_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08083_ (.A1(_06179_),
    .A2(_00370_),
    .B(_00982_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08084_ (.A1(_00984_),
    .A2(_00985_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08085_ (.A1(_05398_),
    .A2(_00376_),
    .B1(_00373_),
    .B2(_05833_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08086_ (.A1(_00987_),
    .A2(_00982_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08087_ (.A1(net58),
    .A2(_06308_),
    .A3(_00355_),
    .A4(net152),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08088_ (.A1(_06308_),
    .A2(_00355_),
    .B1(net152),
    .B2(net58),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08089_ (.I(_00990_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08090_ (.A1(_00991_),
    .A2(_00989_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08091_ (.A1(net73),
    .A2(_05864_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08092_ (.A1(net60),
    .A2(_05833_),
    .B1(_05398_),
    .B2(net61),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08093_ (.A1(net61),
    .A2(net60),
    .A3(_05833_),
    .A4(_05398_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08094_ (.A1(_00993_),
    .A2(_00994_),
    .B(_00995_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08095_ (.A1(_00357_),
    .A2(_06179_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08096_ (.A1(_00363_),
    .A2(_05864_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08097_ (.A1(net61),
    .A2(_05833_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08098_ (.A1(_00997_),
    .A2(_00998_),
    .A3(_00999_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08099_ (.A1(_00996_),
    .A2(_01000_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08100_ (.A1(_00996_),
    .A2(_01000_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08101_ (.A1(_00992_),
    .A2(_01001_),
    .B(_01002_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08102_ (.A1(_00355_),
    .A2(net152),
    .B1(net155),
    .B2(net58),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08103_ (.A1(net58),
    .A2(_00355_),
    .A3(net152),
    .A4(net155),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08104_ (.A1(_01004_),
    .A2(_01005_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08105_ (.A1(net60),
    .A2(_05864_),
    .B1(_05833_),
    .B2(net61),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08106_ (.A1(net61),
    .A2(net60),
    .A3(_05864_),
    .A4(_05833_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08107_ (.A1(_00997_),
    .A2(_01007_),
    .B(_01008_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08108_ (.A1(net158),
    .A2(_05864_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08109_ (.A1(_00363_),
    .A2(_06179_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08110_ (.A1(net73),
    .A2(_06308_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08111_ (.A1(_01010_),
    .A2(_01011_),
    .A3(_01012_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08112_ (.A1(_01009_),
    .A2(_01013_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08113_ (.A1(_01006_),
    .A2(_01014_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08114_ (.A1(_01003_),
    .A2(_01015_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08115_ (.A1(_01003_),
    .A2(_01015_),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08116_ (.A1(_00989_),
    .A2(_01016_),
    .B(_01017_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08117_ (.A1(_01009_),
    .A2(_01013_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08118_ (.A1(_01006_),
    .A2(_01014_),
    .B(_01019_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08119_ (.A1(net137),
    .A2(_06598_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08120_ (.A1(_00355_),
    .A2(net155),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08121_ (.A1(_01021_),
    .A2(_01022_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08122_ (.A1(_01021_),
    .A2(_01022_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08123_ (.A1(_01023_),
    .A2(_01024_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08124_ (.A1(net142),
    .A2(_06179_),
    .B1(_05864_),
    .B2(net61),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08125_ (.A1(net61),
    .A2(net142),
    .A3(_06179_),
    .A4(_05864_),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08126_ (.A1(_01012_),
    .A2(_01026_),
    .B(_01027_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08127_ (.A1(_00363_),
    .A2(_06308_),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08128_ (.A1(net158),
    .A2(_06179_),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08129_ (.A1(net73),
    .A2(_06416_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08130_ (.A1(_01029_),
    .A2(_01030_),
    .A3(_01031_),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08131_ (.A1(_01028_),
    .A2(_01032_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08132_ (.A1(_01025_),
    .A2(_01033_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08133_ (.A1(_01005_),
    .A2(_01020_),
    .A3(_01034_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08134_ (.A1(_01018_),
    .A2(_01035_),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08135_ (.A1(_01018_),
    .A2(_01035_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08136_ (.A1(_00988_),
    .A2(_01036_),
    .B(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08137_ (.A1(_05864_),
    .A2(_00373_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08138_ (.A1(_05833_),
    .A2(_00376_),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08139_ (.A1(_05398_),
    .A2(_00379_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08140_ (.A1(_01040_),
    .A2(_01041_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08141_ (.A1(_01039_),
    .A2(_01042_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08142_ (.A1(net58),
    .A2(_00355_),
    .A3(net152),
    .A4(net155),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08143_ (.A1(_01020_),
    .A2(_01034_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08144_ (.A1(_01020_),
    .A2(_01034_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08145_ (.A1(_01044_),
    .A2(_01045_),
    .B(_01046_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08146_ (.A1(_01028_),
    .A2(_01032_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08147_ (.A1(_01025_),
    .A2(_01033_),
    .B(_01048_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08148_ (.A1(net137),
    .A2(_06618_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08149_ (.A1(_00355_),
    .A2(_06598_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08150_ (.A1(_01050_),
    .A2(_01051_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08151_ (.A1(_01050_),
    .A2(_01051_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08152_ (.A1(_01052_),
    .A2(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08153_ (.A1(net142),
    .A2(_06308_),
    .B1(_06179_),
    .B2(net92),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08154_ (.A1(net91),
    .A2(net142),
    .A3(_06308_),
    .A4(_06179_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08155_ (.A1(_01031_),
    .A2(_01055_),
    .B(_01056_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08156_ (.A1(_00363_),
    .A2(_06416_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08157_ (.A1(_00367_),
    .A2(_06308_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08158_ (.A1(_01058_),
    .A2(_01059_),
    .A3(_00954_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08159_ (.A1(_01060_),
    .A2(_01057_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08160_ (.A1(_01061_),
    .A2(_01054_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08161_ (.A1(_01062_),
    .A2(_01049_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08162_ (.A1(_01024_),
    .A2(_01063_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08163_ (.A1(_01047_),
    .A2(_01064_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08164_ (.A1(_01043_),
    .A2(_01065_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08165_ (.A1(_01038_),
    .A2(_01066_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08166_ (.A1(_01038_),
    .A2(_01066_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08167_ (.A1(_00986_),
    .A2(_01067_),
    .B(_01068_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08168_ (.A1(_01040_),
    .A2(_01041_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08169_ (.A1(_05864_),
    .A2(_00373_),
    .A3(_01042_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08170_ (.A1(_01070_),
    .A2(_01071_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08171_ (.A1(_06308_),
    .A2(_00370_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08172_ (.A1(_01072_),
    .A2(_01073_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08173_ (.A1(_01047_),
    .A2(_01064_),
    .ZN(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08174_ (.A1(_01043_),
    .A2(_01065_),
    .B(_01075_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08175_ (.A1(_05398_),
    .A2(_00382_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08176_ (.A1(_05864_),
    .A2(_05833_),
    .A3(_00379_),
    .A4(_00376_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08177_ (.A1(_05833_),
    .A2(_00379_),
    .B1(_00376_),
    .B2(_05864_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08178_ (.A1(_01078_),
    .A2(_01079_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08179_ (.A1(_06179_),
    .A2(_00373_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08180_ (.A1(_01080_),
    .A2(_01081_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08181_ (.A1(_01077_),
    .A2(_01082_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08182_ (.A1(_01049_),
    .A2(_01062_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08183_ (.A1(_01024_),
    .A2(_01063_),
    .B(_01084_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08184_ (.A1(_01057_),
    .A2(_01060_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08185_ (.A1(_01054_),
    .A2(_01061_),
    .B(_01086_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08186_ (.A1(_00953_),
    .A2(_00961_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08187_ (.A1(_01087_),
    .A2(_01088_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08188_ (.A1(_01053_),
    .A2(_01089_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08189_ (.A1(_01085_),
    .A2(_01090_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08190_ (.A1(_01083_),
    .A2(_01091_),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08191_ (.A1(_01076_),
    .A2(_01092_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08192_ (.A1(_01074_),
    .A2(_01093_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08193_ (.A1(_01069_),
    .A2(_01094_),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08194_ (.A1(_01095_),
    .A2(_00983_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08195_ (.A1(_05864_),
    .A2(_00370_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08196_ (.A1(_05398_),
    .A2(_00373_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08197_ (.A1(net58),
    .A2(_06308_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08198_ (.A1(_00355_),
    .A2(_06179_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08199_ (.A1(_01099_),
    .A2(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08200_ (.A1(net60),
    .A2(net73),
    .A3(_05833_),
    .A4(_05398_),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08201_ (.A1(net142),
    .A2(_05833_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08202_ (.A1(net91),
    .A2(_05398_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08203_ (.A1(_01103_),
    .A2(_01104_),
    .A3(_00993_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08204_ (.A1(_01102_),
    .A2(_01105_),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08205_ (.A1(_01102_),
    .A2(_01105_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08206_ (.A1(_01101_),
    .A2(_01106_),
    .B(_01107_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08207_ (.A1(_00992_),
    .A2(_01001_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08208_ (.A1(_01108_),
    .A2(_01109_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _08209_ (.A1(_01099_),
    .A2(_01100_),
    .A3(_01110_),
    .B1(_01109_),
    .B2(_01108_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08210_ (.A1(_00989_),
    .A2(_01016_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08211_ (.A1(_01111_),
    .A2(_01112_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08212_ (.A1(_01111_),
    .A2(_01112_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08213_ (.A1(_01098_),
    .A2(_01113_),
    .B(_01114_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08214_ (.A1(_00988_),
    .A2(_01036_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08215_ (.A1(_01115_),
    .A2(_01116_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08216_ (.A1(_01115_),
    .A2(_01116_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08217_ (.A1(_01097_),
    .A2(_01117_),
    .B(_01118_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08218_ (.A1(_01038_),
    .A2(_01066_),
    .A3(_00986_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08219_ (.A1(_01119_),
    .A2(_01120_),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08220_ (.A1(_01111_),
    .A2(_01112_),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08221_ (.A1(_01098_),
    .A2(_01122_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08222_ (.A1(_01102_),
    .A2(_01105_),
    .A3(_01101_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08223_ (.A1(net58),
    .A2(_00355_),
    .A3(_06179_),
    .A4(_05864_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08224_ (.A1(net58),
    .A2(_06179_),
    .B1(_05864_),
    .B2(_00355_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08225_ (.A1(_01125_),
    .A2(_01126_),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08226_ (.A1(net73),
    .A2(_05833_),
    .B1(_05398_),
    .B2(net60),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08227_ (.I(_01128_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08228_ (.A1(_01102_),
    .A2(_01129_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08229_ (.A1(_01127_),
    .A2(_01130_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08230_ (.A1(_01125_),
    .A2(_01131_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08231_ (.A1(_01124_),
    .A2(_01132_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08232_ (.A1(_01099_),
    .A2(_01100_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08233_ (.A1(_01134_),
    .A2(_01110_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08234_ (.A1(_01133_),
    .A2(_01135_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08235_ (.A1(_01098_),
    .A2(_01122_),
    .A3(_01136_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08236_ (.A1(_05833_),
    .A2(_00370_),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08237_ (.A1(_01137_),
    .A2(_01138_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08238_ (.A1(_01123_),
    .A2(_01136_),
    .B(_01139_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08239_ (.A1(_01097_),
    .A2(_01117_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08240_ (.A1(_01140_),
    .A2(_01141_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08241_ (.A1(_01119_),
    .A2(_01120_),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08242_ (.A1(_01121_),
    .A2(_01142_),
    .B(_01143_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08243_ (.A1(_01137_),
    .A2(_01138_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08244_ (.A1(_01133_),
    .A2(_01135_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08245_ (.A1(_01124_),
    .A2(_01132_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08246_ (.A1(_01127_),
    .A2(_01130_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08247_ (.A1(net73),
    .A2(_05398_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08248_ (.A1(_00355_),
    .A2(_05833_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08249_ (.A1(_01149_),
    .A2(_01150_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08250_ (.A1(net58),
    .A2(_05864_),
    .A3(_01151_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08251_ (.A1(_01149_),
    .A2(_01150_),
    .B(_01152_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08252_ (.A1(_01147_),
    .A2(_01148_),
    .A3(_01153_),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08253_ (.A1(_01146_),
    .A2(_01154_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08254_ (.I(_01148_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08255_ (.A1(_00993_),
    .A2(_01156_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08256_ (.A1(net58),
    .A2(_00355_),
    .A3(_05833_),
    .A4(_05398_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08257_ (.A1(net73),
    .A2(_05864_),
    .B(_01148_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08258_ (.A1(_01147_),
    .A2(_01157_),
    .A3(_01158_),
    .A4(_01159_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08259_ (.A1(_01155_),
    .A2(_01160_),
    .B(_05398_),
    .C(_00370_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08260_ (.A1(_01155_),
    .A2(_01160_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08261_ (.A1(_01146_),
    .A2(_01154_),
    .B(_01161_),
    .C(_01162_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08262_ (.A1(_01139_),
    .A2(_01141_),
    .A3(_01145_),
    .A4(_01163_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08263_ (.A1(_01121_),
    .A2(_01142_),
    .B(_01164_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08264_ (.A1(_01096_),
    .A2(_01144_),
    .B(_01165_),
    .ZN(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08265_ (.A1(_01119_),
    .A2(_01120_),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08266_ (.A1(_01096_),
    .A2(_01167_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08267_ (.A1(_01069_),
    .A2(_01094_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08268_ (.A1(_00984_),
    .A2(_01095_),
    .B(_01169_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08269_ (.A1(_06308_),
    .A2(_00370_),
    .A3(_01072_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08270_ (.A1(net68),
    .A2(_01092_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08271_ (.A1(_01074_),
    .A2(_01093_),
    .B(_01172_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08272_ (.A1(_01078_),
    .A2(_01079_),
    .A3(_01081_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08273_ (.A1(_01078_),
    .A2(_01174_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08274_ (.A1(net152),
    .A2(_00370_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08275_ (.A1(_01175_),
    .A2(_01176_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08276_ (.A1(_01175_),
    .A2(_01176_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08277_ (.A1(_01177_),
    .A2(_01178_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08278_ (.A1(_01085_),
    .A2(_01090_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08279_ (.A1(_01083_),
    .A2(_01091_),
    .B(_01180_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08280_ (.A1(_01077_),
    .A2(_01082_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08281_ (.A1(_00933_),
    .A2(_00937_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08282_ (.A1(_01182_),
    .A2(_01183_),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08283_ (.I(_01184_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08284_ (.A1(_01087_),
    .A2(_01088_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08285_ (.A1(_01053_),
    .A2(_01089_),
    .B(_01186_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08286_ (.A1(_00951_),
    .A2(_00965_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08287_ (.A1(_01188_),
    .A2(_01187_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08288_ (.A1(_01185_),
    .A2(_01189_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08289_ (.A1(_01181_),
    .A2(_01190_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08290_ (.A1(_01179_),
    .A2(_01191_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08291_ (.A1(_01173_),
    .A2(_01192_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08292_ (.A1(_01171_),
    .A2(_01193_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08293_ (.A1(_01070_),
    .A2(_01071_),
    .B(_01073_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08294_ (.A1(_01173_),
    .A2(_01192_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08295_ (.A1(_01195_),
    .A2(_01193_),
    .B(_01196_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08296_ (.A1(_01181_),
    .A2(_01190_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08297_ (.A1(_01179_),
    .A2(_01191_),
    .B(_01198_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08298_ (.A1(_01182_),
    .A2(_01183_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08299_ (.A1(_00935_),
    .A2(_00936_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08300_ (.A1(_00935_),
    .A2(_00936_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08301_ (.A1(_00934_),
    .A2(_01201_),
    .B(_01202_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08302_ (.A1(net155),
    .A2(_00370_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08303_ (.A1(_01200_),
    .A2(_01203_),
    .A3(_01204_),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08304_ (.I(_01205_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08305_ (.A1(_01187_),
    .A2(_01188_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08306_ (.A1(_01185_),
    .A2(_01189_),
    .B(_01207_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08307_ (.A1(_00948_),
    .A2(_00969_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08308_ (.A1(_01208_),
    .A2(_01209_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08309_ (.A1(_01206_),
    .A2(_01210_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08310_ (.A1(_01177_),
    .A2(_01199_),
    .A3(_01211_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _08311_ (.A1(_01170_),
    .A2(_01194_),
    .B1(_01197_),
    .B2(_01212_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08312_ (.A1(_01166_),
    .A2(_01168_),
    .B(_01213_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08313_ (.A1(_00945_),
    .A2(_00978_),
    .Z(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08314_ (.A1(_01182_),
    .A2(_01183_),
    .B(_01203_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08315_ (.A1(_01182_),
    .A2(_01183_),
    .A3(_01203_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08316_ (.A1(_01216_),
    .A2(_01204_),
    .B(_01217_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08317_ (.I(_01218_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08318_ (.A1(_01208_),
    .A2(_01209_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08319_ (.A1(_01206_),
    .A2(_01210_),
    .B(_01220_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08320_ (.A1(_00947_),
    .A2(_00973_),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _08321_ (.A1(_01222_),
    .A2(_01221_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08322_ (.A1(_01221_),
    .A2(_01222_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08323_ (.A1(_01219_),
    .A2(_01223_),
    .B(_01224_),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08324_ (.A1(_01199_),
    .A2(_01211_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08325_ (.A1(_01199_),
    .A2(_01211_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08326_ (.A1(_01177_),
    .A2(_01226_),
    .B(_01227_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08327_ (.A1(_01219_),
    .A2(_01223_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08328_ (.A1(_01215_),
    .A2(_01225_),
    .B1(_01228_),
    .B2(_01229_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08329_ (.A1(_01173_),
    .A2(_01192_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08330_ (.A1(_01173_),
    .A2(_01192_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08331_ (.A1(_01171_),
    .A2(_01231_),
    .B(_01232_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08332_ (.A1(_01175_),
    .A2(_01176_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _08333_ (.A1(_01234_),
    .A2(_01199_),
    .A3(_01211_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08334_ (.A1(_01195_),
    .A2(_01193_),
    .B(_01235_),
    .C(_01196_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _08335_ (.A1(_01195_),
    .A2(_01173_),
    .A3(_01192_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08336_ (.A1(_00984_),
    .A2(net71),
    .B(_01237_),
    .C(_01169_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08337_ (.A1(_01236_),
    .A2(_01238_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08338_ (.A1(_01233_),
    .A2(_01235_),
    .B(_01239_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08339_ (.A1(_01215_),
    .A2(_01225_),
    .B1(_01228_),
    .B2(_01229_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08340_ (.A1(_01215_),
    .A2(_01225_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08341_ (.A1(_01241_),
    .A2(_01242_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08342_ (.A1(_01214_),
    .A2(_01230_),
    .A3(_01240_),
    .B(_01243_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08343_ (.A1(_00981_),
    .A2(_01244_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08344_ (.A1(_00981_),
    .A2(_01244_),
    .B(_05182_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _08345_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[0] ),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08346_ (.A1(_05280_),
    .A2(_01247_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08347_ (.A1(_01245_),
    .A2(_01246_),
    .B(_01248_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _08348_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[1] ),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08349_ (.A1(_00870_),
    .A2(_00873_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08350_ (.A1(_00874_),
    .A2(_00875_),
    .B(_01250_),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08351_ (.A1(_00878_),
    .A2(_00926_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08352_ (.A1(_00876_),
    .A2(_00927_),
    .B(_01252_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08353_ (.A1(_00880_),
    .A2(_00906_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08354_ (.A1(_00907_),
    .A2(_00925_),
    .B(_01254_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08355_ (.I(_00916_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08356_ (.A1(_00912_),
    .A2(_01256_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08357_ (.A1(_00917_),
    .A2(_00922_),
    .B(_01257_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08358_ (.A1(_00858_),
    .A2(_00881_),
    .B(_00885_),
    .C(_00886_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08359_ (.A1(_00914_),
    .A2(_00915_),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08360_ (.A1(_00914_),
    .A2(_00915_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08361_ (.A1(_00913_),
    .A2(_01260_),
    .B(_01261_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08362_ (.A1(_06523_),
    .A2(_00382_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08363_ (.A1(_06308_),
    .A2(_00388_),
    .ZN(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08364_ (.A1(net153),
    .A2(_00385_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08365_ (.A1(_01263_),
    .A2(_01264_),
    .A3(_01265_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08366_ (.A1(_06627_),
    .A2(_00373_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08367_ (.A1(_06598_),
    .A2(_00379_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08368_ (.A1(_06618_),
    .A2(_00376_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08369_ (.A1(_01268_),
    .A2(_01269_),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08370_ (.A1(_01267_),
    .A2(_01270_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08371_ (.A1(_01262_),
    .A2(_01266_),
    .A3(_01271_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08372_ (.A1(_01259_),
    .A2(_01272_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08373_ (.A1(_01258_),
    .A2(_01273_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08374_ (.A1(_00890_),
    .A2(_00904_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08375_ (.A1(_00888_),
    .A2(_00905_),
    .B(_01275_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08376_ (.A1(_00893_),
    .A2(_00897_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08377_ (.A1(_00898_),
    .A2(_00903_),
    .B(_01277_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08378_ (.A1(net143),
    .A2(_06637_),
    .B1(_06633_),
    .B2(net91),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08379_ (.A1(net91),
    .A2(net143),
    .A3(_06637_),
    .A4(_06633_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08380_ (.A1(_00894_),
    .A2(_01279_),
    .B(_01280_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08381_ (.A1(_06649_),
    .A2(_00357_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08382_ (.A1(_00367_),
    .A2(_06637_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08383_ (.A1(_06642_),
    .A2(_00363_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08384_ (.A1(_01282_),
    .A2(_01283_),
    .A3(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08385_ (.A1(_01285_),
    .A2(_01281_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08386_ (.A1(_06654_),
    .A2(_00355_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08387_ (.A1(_00352_),
    .A2(_06659_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08388_ (.A1(net96),
    .A2(_06179_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08389_ (.A1(_01287_),
    .A2(_01288_),
    .A3(_01289_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08390_ (.A1(_01286_),
    .A2(_01290_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08391_ (.A1(_00899_),
    .A2(_00900_),
    .A3(_00901_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08392_ (.A1(_00900_),
    .A2(_01292_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08393_ (.A1(_00398_),
    .A2(_05833_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08394_ (.A1(_05864_),
    .A2(_00394_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08395_ (.A1(_01293_),
    .A2(_01294_),
    .A3(_01295_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08396_ (.A1(_00885_),
    .A2(_01296_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08397_ (.A1(_01278_),
    .A2(_01291_),
    .A3(_01297_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08398_ (.A1(_01276_),
    .A2(_01298_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08399_ (.A1(_01274_),
    .A2(_01299_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08400_ (.A1(_06633_),
    .A2(_00370_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08401_ (.A1(_00394_),
    .A2(_05398_),
    .A3(_00844_),
    .A4(_00923_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08402_ (.A1(_00909_),
    .A2(_00924_),
    .B(_01302_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08403_ (.A1(_00919_),
    .A2(_00920_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08404_ (.A1(_00918_),
    .A2(_00921_),
    .B(_01304_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08405_ (.A1(_01303_),
    .A2(_01305_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08406_ (.A1(_01301_),
    .A2(_01306_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08407_ (.A1(_01255_),
    .A2(_01300_),
    .A3(_01307_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08408_ (.A1(_01253_),
    .A2(_01308_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08409_ (.A1(_01309_),
    .A2(_01251_),
    .Z(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08410_ (.A1(_00869_),
    .A2(_00928_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08411_ (.A1(_00869_),
    .A2(_00928_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08412_ (.A1(_00768_),
    .A2(_01311_),
    .B(_01312_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08413_ (.A1(_01310_),
    .A2(_01313_),
    .Z(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08414_ (.A1(_00930_),
    .A2(_00980_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08415_ (.A1(_00981_),
    .A2(_01244_),
    .B(_01315_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _08416_ (.A1(_01314_),
    .A2(_01316_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08417_ (.A1(_00418_),
    .A2(_01317_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08418_ (.I0(_01249_),
    .I1(_01318_),
    .S(_00395_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08419_ (.I(_01319_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08420_ (.A1(_00418_),
    .A2(_01317_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08421_ (.A1(_00767_),
    .A2(_00929_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _08422_ (.A1(_01312_),
    .A2(_01321_),
    .A3(_01310_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _08423_ (.A1(_00980_),
    .A2(_00930_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08424_ (.A1(_01323_),
    .A2(_01314_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08425_ (.A1(_01241_),
    .A2(_01242_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08426_ (.I(_01310_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08427_ (.A1(_01326_),
    .A2(_01313_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08428_ (.A1(_01315_),
    .A2(_01322_),
    .B1(_01324_),
    .B2(_01325_),
    .C(_01327_),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08429_ (.A1(_01069_),
    .A2(_01094_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08430_ (.A1(_01069_),
    .A2(_01094_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08431_ (.A1(_00983_),
    .A2(_01329_),
    .B(_01330_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08432_ (.A1(_01331_),
    .A2(_01237_),
    .B1(_01233_),
    .B2(_01235_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _08433_ (.A1(_01096_),
    .A2(_01144_),
    .A3(_01238_),
    .Z(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08434_ (.A1(_01332_),
    .A2(_01333_),
    .B(_01236_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08435_ (.A1(_01236_),
    .A2(_01165_),
    .Z(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08436_ (.A1(_01143_),
    .A2(_01096_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08437_ (.A1(_01213_),
    .A2(_01238_),
    .A3(_01335_),
    .A4(_01336_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08438_ (.A1(_00945_),
    .A2(_00978_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08439_ (.A1(_01221_),
    .A2(_01222_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08440_ (.A1(_01221_),
    .A2(_01222_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08441_ (.A1(_01218_),
    .A2(_01339_),
    .B(_01340_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08442_ (.A1(_01199_),
    .A2(_01211_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08443_ (.A1(_01199_),
    .A2(_01211_),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08444_ (.A1(_01234_),
    .A2(_01342_),
    .B(_01343_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08445_ (.A1(_01218_),
    .A2(_01223_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08446_ (.A1(_01338_),
    .A2(_01341_),
    .B1(_01344_),
    .B2(_01345_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08447_ (.A1(_01346_),
    .A2(_01230_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _08448_ (.A1(_01334_),
    .A2(_01337_),
    .B(_01347_),
    .C(_01324_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08449_ (.A1(_01348_),
    .A2(_01328_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08450_ (.A1(_06633_),
    .A2(_00370_),
    .A3(_01306_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08451_ (.A1(_01303_),
    .A2(_01305_),
    .B(_01350_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08452_ (.A1(_01255_),
    .A2(_01300_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08453_ (.A1(_01255_),
    .A2(_01300_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08454_ (.A1(_01352_),
    .A2(_01307_),
    .B(_01353_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08455_ (.I(_01273_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08456_ (.A1(_01259_),
    .A2(_01272_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08457_ (.A1(_01258_),
    .A2(_01355_),
    .B(_01356_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08458_ (.A1(_01268_),
    .A2(_01269_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08459_ (.A1(_06627_),
    .A2(_00373_),
    .A3(_01270_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08460_ (.A1(_01358_),
    .A2(_01359_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08461_ (.A1(_01357_),
    .A2(_01360_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08462_ (.A1(_06637_),
    .A2(_00370_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08463_ (.A1(_01361_),
    .A2(_01362_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08464_ (.I(_01274_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08465_ (.A1(_01276_),
    .A2(_01298_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08466_ (.A1(_01364_),
    .A2(_01299_),
    .B(_01365_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08467_ (.A1(_01262_),
    .A2(_01266_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08468_ (.A1(_01262_),
    .A2(_01266_),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08469_ (.A1(_01367_),
    .A2(_01271_),
    .B(_01368_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08470_ (.A1(_01294_),
    .A2(_01295_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08471_ (.A1(_01294_),
    .A2(_01295_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08472_ (.A1(_01293_),
    .A2(_01370_),
    .A3(_01371_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08473_ (.A1(_00885_),
    .A2(_01296_),
    .B(_01372_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08474_ (.A1(_06633_),
    .A2(_00373_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08475_ (.A1(_00379_),
    .A2(_06618_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08476_ (.A1(_06627_),
    .A2(_00376_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08477_ (.A1(_01375_),
    .A2(_01376_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08478_ (.A1(_01374_),
    .A2(_01377_),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08479_ (.A1(_01264_),
    .A2(_01265_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08480_ (.A1(_01264_),
    .A2(_01265_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08481_ (.A1(_01263_),
    .A2(_01379_),
    .B(_01380_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08482_ (.A1(_00382_),
    .A2(_06598_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08483_ (.A1(_00388_),
    .A2(_06416_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08484_ (.A1(_00385_),
    .A2(net156),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08485_ (.A1(_01382_),
    .A2(_01383_),
    .A3(_01384_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08486_ (.A1(_01381_),
    .A2(_01385_),
    .Z(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08487_ (.A1(_01378_),
    .A2(_01386_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08488_ (.A1(_01373_),
    .A2(_01387_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08489_ (.A1(_01369_),
    .A2(_01388_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08490_ (.A1(_01278_),
    .A2(_01291_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08491_ (.A1(_01278_),
    .A2(_01291_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08492_ (.A1(_01390_),
    .A2(_01297_),
    .B(_01391_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08493_ (.A1(_01288_),
    .A2(_01289_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08494_ (.A1(_01288_),
    .A2(_01289_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08495_ (.A1(_01287_),
    .A2(_01393_),
    .B(_01394_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08496_ (.A1(_00398_),
    .A2(_05864_),
    .B1(_00394_),
    .B2(_06179_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08497_ (.A1(_06179_),
    .A2(_00398_),
    .A3(_05864_),
    .A4(_00394_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08498_ (.A1(_01396_),
    .A2(_01397_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08499_ (.A1(_01371_),
    .A2(_01395_),
    .A3(_01398_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08500_ (.A1(_01281_),
    .A2(_01285_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08501_ (.A1(net154),
    .A2(_01290_),
    .B(_01400_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08502_ (.A1(_00355_),
    .A2(_06659_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08503_ (.A1(net58),
    .A2(_06664_),
    .A3(net95),
    .A4(_06308_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08504_ (.A1(net137),
    .A2(_06664_),
    .B1(net95),
    .B2(_06308_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08505_ (.A1(_01403_),
    .A2(_01404_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08506_ (.A1(_01402_),
    .A2(_01405_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08507_ (.A1(_06642_),
    .A2(net60),
    .B1(_06637_),
    .B2(net61),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08508_ (.A1(_06642_),
    .A2(net61),
    .A3(net60),
    .A4(_06637_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08509_ (.A1(_01282_),
    .A2(_01407_),
    .B(_01408_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08510_ (.A1(_00357_),
    .A2(_06654_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08511_ (.A1(_06642_),
    .A2(net91),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08512_ (.A1(net60),
    .A2(_06649_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08513_ (.A1(_01410_),
    .A2(_01411_),
    .A3(_01412_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08514_ (.A1(_01409_),
    .A2(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08515_ (.A1(_01406_),
    .A2(_01414_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08516_ (.A1(_01399_),
    .A2(_01401_),
    .A3(_01415_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08517_ (.A1(_01392_),
    .A2(_01416_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08518_ (.A1(_01389_),
    .A2(_01417_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08519_ (.A1(_01366_),
    .A2(_01418_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08520_ (.A1(_01363_),
    .A2(_01419_),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08521_ (.A1(_01354_),
    .A2(_01420_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08522_ (.A1(_01351_),
    .A2(_01421_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08523_ (.A1(_01253_),
    .A2(_01308_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08524_ (.A1(_01251_),
    .A2(_01309_),
    .B(_01423_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08525_ (.A1(_01422_),
    .A2(_01424_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _08526_ (.A1(_00424_),
    .A2(_01349_),
    .A3(_01425_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08527_ (.A1(_01320_),
    .A2(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08528_ (.A1(_01320_),
    .A2(_01426_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08529_ (.A1(_05182_),
    .A2(_01428_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _08530_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[2] ),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08531_ (.A1(_05280_),
    .A2(_01430_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08532_ (.A1(_01427_),
    .A2(_01429_),
    .B(_01431_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08533_ (.I(_01425_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08534_ (.A1(net56),
    .A2(_01348_),
    .B(_01432_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08535_ (.A1(_01349_),
    .A2(_01425_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_4 _08536_ (.A1(_00424_),
    .A2(_01433_),
    .A3(_01434_),
    .B1(_01426_),
    .B2(_01317_),
    .B3(_00418_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08537_ (.A1(_01354_),
    .A2(_01420_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08538_ (.A1(_01351_),
    .A2(_01421_),
    .B(_01436_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08539_ (.A1(_01358_),
    .A2(_01359_),
    .B(_01357_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08540_ (.A1(_01361_),
    .A2(_01362_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08541_ (.A1(_01438_),
    .A2(_01439_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08542_ (.A1(_01366_),
    .A2(_01418_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08543_ (.A1(_01363_),
    .A2(_01419_),
    .B(_01441_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08544_ (.A1(_01373_),
    .A2(_01387_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08545_ (.A1(_01369_),
    .A2(_01388_),
    .B(_01443_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08546_ (.A1(_01375_),
    .A2(_01376_),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08547_ (.A1(_06633_),
    .A2(_00373_),
    .A3(_01377_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08548_ (.A1(_01445_),
    .A2(_01446_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08549_ (.A1(_01447_),
    .A2(_01444_),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08550_ (.A1(_06642_),
    .A2(_00370_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08551_ (.A1(_01448_),
    .A2(_01449_),
    .Z(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08552_ (.A1(_01392_),
    .A2(_01416_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08553_ (.A1(_01389_),
    .A2(_01417_),
    .B(_01451_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08554_ (.I(_01385_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08555_ (.A1(_01381_),
    .A2(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08556_ (.A1(_01378_),
    .A2(_01386_),
    .B(_01454_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08557_ (.A1(_01395_),
    .A2(_01398_),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08558_ (.A1(_01395_),
    .A2(_01398_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08559_ (.A1(_01371_),
    .A2(_01456_),
    .B(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08560_ (.A1(_06637_),
    .A2(_00373_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08561_ (.A1(_06627_),
    .A2(_00379_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08562_ (.A1(_06633_),
    .A2(_00376_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08563_ (.A1(_01460_),
    .A2(_01461_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08564_ (.A1(_01459_),
    .A2(_01462_),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08565_ (.A1(_01383_),
    .A2(_01384_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08566_ (.A1(_01383_),
    .A2(_01384_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08567_ (.A1(_01382_),
    .A2(_01464_),
    .B(_01465_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08568_ (.A1(_00382_),
    .A2(_06618_),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08569_ (.A1(_00388_),
    .A2(_06523_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08570_ (.A1(_00385_),
    .A2(_06598_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08571_ (.A1(_01467_),
    .A2(_01468_),
    .A3(_01469_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08572_ (.A1(_01466_),
    .A2(_01470_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08573_ (.A1(_01463_),
    .A2(_01471_),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08574_ (.A1(_01458_),
    .A2(_01472_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08575_ (.A1(_01455_),
    .A2(_01473_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08576_ (.A1(_01401_),
    .A2(_01415_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08577_ (.A1(_01401_),
    .A2(_01415_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08578_ (.A1(_01399_),
    .A2(_01475_),
    .B(_01476_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08579_ (.A1(net58),
    .A2(_06664_),
    .A3(net95),
    .A4(_06308_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08580_ (.A1(_01402_),
    .A2(_01404_),
    .B(_01478_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08581_ (.A1(_06179_),
    .A2(_00398_),
    .B1(_00394_),
    .B2(_06308_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08582_ (.A1(_06308_),
    .A2(_06179_),
    .A3(_00398_),
    .A4(_00394_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08583_ (.A1(_01480_),
    .A2(_01481_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08584_ (.A1(_01479_),
    .A2(_01482_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08585_ (.A1(_01397_),
    .A2(_01483_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08586_ (.A1(_01409_),
    .A2(_01413_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08587_ (.A1(_01406_),
    .A2(_01414_),
    .B(_01485_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08588_ (.A1(_06642_),
    .A2(net61),
    .B1(net60),
    .B2(_06649_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08589_ (.A1(_06642_),
    .A2(net61),
    .A3(net60),
    .A4(_06649_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08590_ (.A1(_01410_),
    .A2(_01487_),
    .B(_01488_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08591_ (.A1(net73),
    .A2(_06659_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08592_ (.A1(net91),
    .A2(_06649_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08593_ (.A1(net60),
    .A2(_06654_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08594_ (.A1(_01490_),
    .A2(_01491_),
    .A3(_01492_),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08595_ (.A1(_01489_),
    .A2(_01493_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08596_ (.A1(net58),
    .A2(net95),
    .A3(net152),
    .A4(_06672_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08597_ (.A1(net97),
    .A2(net153),
    .B1(_06672_),
    .B2(net137),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08598_ (.A1(_01495_),
    .A2(_01496_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08599_ (.A1(_06664_),
    .A2(_00355_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08600_ (.A1(_01497_),
    .A2(_01498_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08601_ (.A1(_01494_),
    .A2(_01499_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08602_ (.A1(_01484_),
    .A2(_01486_),
    .A3(_01500_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08603_ (.A1(_01477_),
    .A2(_01501_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08604_ (.A1(_01474_),
    .A2(_01502_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08605_ (.A1(_01450_),
    .A2(_01452_),
    .A3(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08606_ (.A1(_01442_),
    .A2(_01504_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _08607_ (.A1(_01440_),
    .A2(_01505_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08608_ (.A1(_01437_),
    .A2(_01506_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08609_ (.I(_01507_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08610_ (.A1(_01422_),
    .A2(_01424_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08611_ (.I(_01509_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _08612_ (.A1(_01314_),
    .A2(_01323_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08613_ (.A1(_01315_),
    .A2(_01322_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _08614_ (.A1(_01326_),
    .A2(_01313_),
    .B1(_01511_),
    .B2(_01243_),
    .C(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08615_ (.A1(_01096_),
    .A2(_01144_),
    .A3(_01238_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08616_ (.A1(_01233_),
    .A2(_01235_),
    .B1(_01213_),
    .B2(_01514_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _08617_ (.A1(_01213_),
    .A2(_01238_),
    .A3(_01335_),
    .A4(_01336_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08618_ (.A1(_01346_),
    .A2(_01230_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08619_ (.A1(_01515_),
    .A2(_01516_),
    .B(_01517_),
    .C(_01511_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08620_ (.A1(_01513_),
    .A2(_01518_),
    .B(_01425_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08621_ (.A1(_01510_),
    .A2(_01519_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _08622_ (.A1(_00428_),
    .A2(_01508_),
    .A3(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08623_ (.A1(_01435_),
    .A2(_01521_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08624_ (.A1(_01435_),
    .A2(_01521_),
    .B(_05182_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _08625_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[3] ),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08626_ (.A1(_05280_),
    .A2(_01524_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08627_ (.A1(_01522_),
    .A2(_01523_),
    .B(_01525_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08628_ (.A1(_01510_),
    .A2(_01519_),
    .B(_01508_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08629_ (.A1(_01509_),
    .A2(_01433_),
    .A3(_01507_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08630_ (.A1(_00428_),
    .A2(_01526_),
    .A3(_01527_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08631_ (.A1(_01435_),
    .A2(_01521_),
    .B(_01528_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08632_ (.A1(_01437_),
    .A2(_01506_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08633_ (.A1(_01422_),
    .A2(_01424_),
    .B1(_01437_),
    .B2(_01506_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08634_ (.A1(_01530_),
    .A2(_01531_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08635_ (.I(_01532_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08636_ (.A1(_01328_),
    .A2(_01348_),
    .B(_01432_),
    .C(_01508_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08637_ (.A1(_01445_),
    .A2(_01446_),
    .B(_01444_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08638_ (.A1(_01448_),
    .A2(_01449_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08639_ (.A1(_01535_),
    .A2(_01536_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08640_ (.A1(_01452_),
    .A2(_01503_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08641_ (.A1(_01452_),
    .A2(_01503_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08642_ (.A1(_01450_),
    .A2(_01538_),
    .B(_01539_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08643_ (.A1(_01458_),
    .A2(_01472_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08644_ (.A1(_01455_),
    .A2(_01473_),
    .B(_01541_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08645_ (.A1(_01460_),
    .A2(_01461_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08646_ (.A1(_06637_),
    .A2(_00373_),
    .A3(_01462_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08647_ (.A1(_01543_),
    .A2(_01544_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08648_ (.A1(_01542_),
    .A2(_01545_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08649_ (.A1(_06649_),
    .A2(_00370_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08650_ (.A1(_01546_),
    .A2(_01547_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08651_ (.A1(_01477_),
    .A2(_01501_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08652_ (.A1(_01474_),
    .A2(_01502_),
    .B(_01549_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08653_ (.A1(_01466_),
    .A2(_01470_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08654_ (.A1(_01463_),
    .A2(_01471_),
    .B(_01551_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08655_ (.A1(_01479_),
    .A2(_01482_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08656_ (.A1(_01397_),
    .A2(_01483_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08657_ (.A1(_01553_),
    .A2(_01554_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08658_ (.A1(_06642_),
    .A2(_00373_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08659_ (.A1(_06633_),
    .A2(_00379_),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08660_ (.A1(_06637_),
    .A2(_00376_),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08661_ (.A1(_01557_),
    .A2(_01558_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08662_ (.A1(_01556_),
    .A2(_01559_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08663_ (.A1(_01468_),
    .A2(_01469_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08664_ (.A1(_01468_),
    .A2(_01469_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08665_ (.A1(_01467_),
    .A2(_01561_),
    .B(_01562_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08666_ (.A1(_06627_),
    .A2(_00382_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08667_ (.A1(_00388_),
    .A2(_06598_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08668_ (.A1(_00385_),
    .A2(_06618_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08669_ (.A1(_01564_),
    .A2(_01565_),
    .A3(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08670_ (.A1(_01563_),
    .A2(_01567_),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08671_ (.A1(_01560_),
    .A2(_01568_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08672_ (.A1(_01555_),
    .A2(_01569_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08673_ (.A1(_01552_),
    .A2(_01570_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08674_ (.A1(_01486_),
    .A2(_01500_),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08675_ (.A1(_01486_),
    .A2(_01500_),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08676_ (.A1(_01484_),
    .A2(_01572_),
    .B(_01573_),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08677_ (.A1(net137),
    .A2(net96),
    .A3(net152),
    .A4(_06672_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08678_ (.A1(_01496_),
    .A2(_01498_),
    .B(_01575_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08679_ (.A1(_06308_),
    .A2(_00398_),
    .B1(_00394_),
    .B2(net152),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08680_ (.A1(_06308_),
    .A2(_00398_),
    .A3(_00394_),
    .A4(net153),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08681_ (.A1(_01577_),
    .A2(_01578_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08682_ (.A1(_01579_),
    .A2(_01576_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08683_ (.A1(_01481_),
    .A2(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08684_ (.A1(_01489_),
    .A2(_01493_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08685_ (.A1(_01494_),
    .A2(_01499_),
    .B(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08686_ (.A1(_00355_),
    .A2(_06672_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08687_ (.A1(net137),
    .A2(_06674_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08688_ (.A1(net95),
    .A2(net155),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08689_ (.A1(_01584_),
    .A2(_01585_),
    .A3(_01586_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08690_ (.A1(net61),
    .A2(_06649_),
    .B1(_06654_),
    .B2(net60),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08691_ (.A1(net61),
    .A2(net60),
    .A3(_06649_),
    .A4(_06654_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08692_ (.A1(_01490_),
    .A2(_01588_),
    .B(_01589_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08693_ (.A1(net73),
    .A2(_06664_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08694_ (.A1(net91),
    .A2(_06654_),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08695_ (.A1(net60),
    .A2(_06659_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08696_ (.A1(_01591_),
    .A2(_01592_),
    .A3(_01593_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08697_ (.A1(_01590_),
    .A2(_01594_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08698_ (.A1(_01587_),
    .A2(_01595_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08699_ (.A1(_01581_),
    .A2(_01583_),
    .A3(_01596_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08700_ (.A1(_01574_),
    .A2(_01597_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08701_ (.A1(_01571_),
    .A2(_01598_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08702_ (.A1(_01548_),
    .A2(_01550_),
    .A3(_01599_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08703_ (.A1(_01540_),
    .A2(_01600_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08704_ (.A1(_01537_),
    .A2(_01601_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08705_ (.A1(_01442_),
    .A2(_01504_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08706_ (.A1(_01440_),
    .A2(_01505_),
    .B(_01603_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08707_ (.A1(_01602_),
    .A2(_01604_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08708_ (.A1(_01533_),
    .A2(_01534_),
    .B(_01605_),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08709_ (.A1(_01605_),
    .A2(_01533_),
    .A3(_01534_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08710_ (.A1(_01606_),
    .A2(_01607_),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08711_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-22] ),
    .A2(_01529_),
    .A3(_01608_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _08712_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[4] ),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08713_ (.A1(_05280_),
    .A2(_01610_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08714_ (.A1(_06059_),
    .A2(_01609_),
    .B(_01611_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08715_ (.A1(_01602_),
    .A2(_01604_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08716_ (.I(_01612_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08717_ (.A1(_01613_),
    .A2(_01606_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08718_ (.A1(_01540_),
    .A2(_01600_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08719_ (.A1(_01537_),
    .A2(_01601_),
    .B(_01615_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08720_ (.A1(_01543_),
    .A2(_01544_),
    .B(_01542_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08721_ (.A1(_01546_),
    .A2(_01547_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08722_ (.A1(_01617_),
    .A2(_01618_),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08723_ (.A1(_01550_),
    .A2(_01599_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08724_ (.A1(_01550_),
    .A2(_01599_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08725_ (.A1(_01548_),
    .A2(_01620_),
    .B(_01621_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08726_ (.A1(_01555_),
    .A2(_01569_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08727_ (.A1(_01552_),
    .A2(_01570_),
    .B(_01623_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08728_ (.A1(_01557_),
    .A2(_01558_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08729_ (.A1(_06642_),
    .A2(_00373_),
    .A3(_01559_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08730_ (.A1(_01625_),
    .A2(_01626_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08731_ (.A1(_01624_),
    .A2(_01627_),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08732_ (.A1(_06654_),
    .A2(_00370_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08733_ (.A1(_01628_),
    .A2(_01629_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08734_ (.A1(_01574_),
    .A2(_01597_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08735_ (.A1(_01571_),
    .A2(_01598_),
    .B(_01631_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08736_ (.A1(_01563_),
    .A2(_01567_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08737_ (.A1(_01560_),
    .A2(_01568_),
    .B(_01633_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08738_ (.A1(_01576_),
    .A2(_01579_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08739_ (.A1(_01481_),
    .A2(_01580_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08740_ (.A1(_01635_),
    .A2(_01636_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08741_ (.A1(_06649_),
    .A2(_00373_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08742_ (.A1(_06637_),
    .A2(_00379_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08743_ (.A1(_06642_),
    .A2(_00376_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08744_ (.A1(_01639_),
    .A2(_01640_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08745_ (.A1(_01638_),
    .A2(_01641_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08746_ (.A1(_01565_),
    .A2(_01566_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08747_ (.A1(_01565_),
    .A2(_01566_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08748_ (.A1(_01564_),
    .A2(_01643_),
    .B(_01644_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08749_ (.A1(_06633_),
    .A2(_00382_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08750_ (.A1(_00388_),
    .A2(_06618_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08751_ (.A1(_06627_),
    .A2(_00385_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08752_ (.A1(_01646_),
    .A2(_01647_),
    .A3(_01648_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08753_ (.A1(_01645_),
    .A2(_01649_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08754_ (.A1(_01642_),
    .A2(_01650_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08755_ (.A1(_01637_),
    .A2(_01651_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08756_ (.A1(_01634_),
    .A2(_01652_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08757_ (.A1(_01583_),
    .A2(_01596_),
    .ZN(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08758_ (.A1(_01583_),
    .A2(_01596_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08759_ (.A1(_01581_),
    .A2(_01654_),
    .B(_01655_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08760_ (.A1(net95),
    .A2(net155),
    .B1(_06674_),
    .B2(net137),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08761_ (.A1(net58),
    .A2(net95),
    .A3(net155),
    .A4(_06674_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08762_ (.A1(_01584_),
    .A2(_01657_),
    .B(_01658_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08763_ (.A1(_00398_),
    .A2(net153),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08764_ (.A1(_00394_),
    .A2(net156),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08765_ (.A1(_01660_),
    .A2(_01661_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08766_ (.A1(_01659_),
    .A2(_01662_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08767_ (.A1(_01578_),
    .A2(_01663_),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08768_ (.A1(_01590_),
    .A2(_01594_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08769_ (.A1(_01587_),
    .A2(_01595_),
    .B(_01665_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08770_ (.A1(_00355_),
    .A2(_06674_),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08771_ (.A1(net137),
    .A2(_06679_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08772_ (.A1(net95),
    .A2(_06598_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08773_ (.A1(_01667_),
    .A2(_01668_),
    .A3(_01669_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08774_ (.A1(net61),
    .A2(_06654_),
    .B1(_06659_),
    .B2(net60),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08775_ (.A1(net61),
    .A2(net60),
    .A3(_06654_),
    .A4(_06659_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08776_ (.A1(_01591_),
    .A2(_01671_),
    .B(_01672_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08777_ (.A1(net73),
    .A2(_06672_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08778_ (.A1(net91),
    .A2(_06659_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08779_ (.A1(net60),
    .A2(_06664_),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08780_ (.A1(_01674_),
    .A2(_01675_),
    .A3(_01676_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08781_ (.A1(_01673_),
    .A2(_01677_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08782_ (.A1(_01670_),
    .A2(_01678_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08783_ (.A1(_01664_),
    .A2(_01666_),
    .A3(_01679_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08784_ (.A1(_01656_),
    .A2(_01680_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08785_ (.A1(_01653_),
    .A2(_01681_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08786_ (.A1(_01632_),
    .A2(_01682_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08787_ (.A1(_01630_),
    .A2(_01683_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08788_ (.A1(_01619_),
    .A2(_01622_),
    .A3(_01684_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08789_ (.I(_01685_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08790_ (.A1(_01616_),
    .A2(_01686_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _08791_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-21] ),
    .A2(_01614_),
    .A3(_01687_),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08792_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-22] ),
    .A2(_01608_),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08793_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-22] ),
    .A2(_01608_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08794_ (.A1(_01529_),
    .A2(_01689_),
    .B(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08795_ (.A1(_01688_),
    .A2(_01691_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _08796_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[5] ),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08797_ (.A1(_05280_),
    .A2(_01693_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08798_ (.A1(_06059_),
    .A2(_01692_),
    .B(_01694_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08799_ (.A1(_01530_),
    .A2(_01605_),
    .A3(_01531_),
    .A4(_01687_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08800_ (.A1(_01616_),
    .A2(_01686_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08801_ (.A1(_01616_),
    .A2(_01686_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08802_ (.A1(_01612_),
    .A2(_01696_),
    .B(_01697_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08803_ (.A1(_01695_),
    .A2(_01698_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08804_ (.A1(_01425_),
    .A2(_01507_),
    .A3(_01605_),
    .A4(_01687_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08805_ (.A1(net56),
    .A2(_01348_),
    .B(_01700_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08806_ (.A1(_01625_),
    .A2(_01626_),
    .B(_01624_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08807_ (.A1(_01628_),
    .A2(_01629_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08808_ (.A1(_01702_),
    .A2(_01703_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08809_ (.A1(_01632_),
    .A2(_01682_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08810_ (.A1(_01630_),
    .A2(_01683_),
    .B(_01705_),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08811_ (.A1(_01637_),
    .A2(_01651_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08812_ (.A1(_01634_),
    .A2(_01652_),
    .B(_01707_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08813_ (.A1(_01639_),
    .A2(_01640_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08814_ (.A1(_06649_),
    .A2(_00373_),
    .A3(_01641_),
    .ZN(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08815_ (.A1(_01709_),
    .A2(_01710_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08816_ (.A1(_01708_),
    .A2(_01711_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08817_ (.A1(_06659_),
    .A2(_00370_),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08818_ (.A1(_01712_),
    .A2(_01713_),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08819_ (.A1(_01656_),
    .A2(_01680_),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08820_ (.A1(_01653_),
    .A2(_01681_),
    .B(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08821_ (.A1(_01645_),
    .A2(_01649_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08822_ (.A1(_01642_),
    .A2(_01650_),
    .B(_01717_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08823_ (.A1(_01659_),
    .A2(_01662_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08824_ (.A1(_01578_),
    .A2(_01663_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08825_ (.A1(_01719_),
    .A2(_01720_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08826_ (.A1(_06654_),
    .A2(_00373_),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08827_ (.A1(_06642_),
    .A2(_00379_),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08828_ (.A1(_06649_),
    .A2(_00376_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08829_ (.A1(_01723_),
    .A2(_01724_),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08830_ (.A1(_01722_),
    .A2(_01725_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08831_ (.A1(_01647_),
    .A2(_01648_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08832_ (.A1(_01647_),
    .A2(_01648_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08833_ (.A1(_01646_),
    .A2(_01727_),
    .B(_01728_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08834_ (.A1(_06637_),
    .A2(_00382_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08835_ (.A1(_06627_),
    .A2(_00388_),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08836_ (.A1(_06633_),
    .A2(_00385_),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08837_ (.A1(_01730_),
    .A2(_01731_),
    .A3(_01732_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08838_ (.A1(_01729_),
    .A2(_01733_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08839_ (.A1(_01726_),
    .A2(_01734_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08840_ (.A1(_01721_),
    .A2(_01735_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08841_ (.A1(_01718_),
    .A2(_01736_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08842_ (.A1(_01666_),
    .A2(_01679_),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08843_ (.A1(_01666_),
    .A2(_01679_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08844_ (.A1(_01664_),
    .A2(_01738_),
    .B(_01739_),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08845_ (.A1(_01660_),
    .A2(_01661_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08846_ (.A1(_01668_),
    .A2(_01669_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08847_ (.A1(_01668_),
    .A2(_01669_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08848_ (.A1(_01667_),
    .A2(_01742_),
    .B(_01743_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08849_ (.A1(_00398_),
    .A2(net155),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08850_ (.A1(_00394_),
    .A2(_06598_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08851_ (.A1(_01745_),
    .A2(_01746_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08852_ (.A1(_01741_),
    .A2(_01744_),
    .A3(_01747_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08853_ (.A1(_01673_),
    .A2(_01677_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08854_ (.A1(_01670_),
    .A2(_01678_),
    .B(_01749_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08855_ (.A1(_00355_),
    .A2(_06679_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08856_ (.A1(net138),
    .A2(_06685_),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08857_ (.A1(net96),
    .A2(_06618_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08858_ (.A1(_01751_),
    .A2(_01752_),
    .A3(_01753_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08859_ (.A1(net60),
    .A2(_06664_),
    .B1(_06659_),
    .B2(net61),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08860_ (.A1(net61),
    .A2(net60),
    .A3(_06664_),
    .A4(_06659_),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08861_ (.A1(_01674_),
    .A2(_01755_),
    .B(_01756_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08862_ (.A1(_00357_),
    .A2(_06674_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08863_ (.A1(net92),
    .A2(_06664_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08864_ (.A1(net60),
    .A2(_06672_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08865_ (.A1(_01758_),
    .A2(_01759_),
    .A3(_01760_),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08866_ (.A1(_01757_),
    .A2(_01761_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08867_ (.A1(_01754_),
    .A2(_01762_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08868_ (.A1(_01750_),
    .A2(_01763_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08869_ (.A1(_01748_),
    .A2(_01764_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08870_ (.A1(_01740_),
    .A2(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08871_ (.A1(_01737_),
    .A2(_01766_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08872_ (.A1(_01716_),
    .A2(_01767_),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08873_ (.A1(_01714_),
    .A2(_01768_),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08874_ (.A1(_01704_),
    .A2(_01706_),
    .A3(_01769_),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08875_ (.A1(_01622_),
    .A2(_01684_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08876_ (.A1(_01622_),
    .A2(_01684_),
    .ZN(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08877_ (.A1(_01619_),
    .A2(_01771_),
    .B(_01772_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08878_ (.A1(_01770_),
    .A2(_01773_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08879_ (.A1(_01699_),
    .A2(_01701_),
    .B(_01774_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08880_ (.I(_01699_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08881_ (.A1(_01425_),
    .A2(_01507_),
    .A3(_01605_),
    .A4(_01687_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08882_ (.A1(_01513_),
    .A2(_01518_),
    .B(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08883_ (.I(_01774_),
    .ZN(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08884_ (.A1(_01776_),
    .A2(_01778_),
    .A3(_01779_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08885_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-20] ),
    .A2(_01775_),
    .A3(_01780_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08886_ (.A1(_01775_),
    .A2(_01780_),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08887_ (.A1(_00440_),
    .A2(_01782_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08888_ (.A1(_01781_),
    .A2(_01783_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08889_ (.A1(_01613_),
    .A2(_01606_),
    .B(_01687_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08890_ (.A1(_01613_),
    .A2(_01606_),
    .A3(_01687_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08891_ (.A1(_01785_),
    .A2(_01786_),
    .B(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-21] ),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08892_ (.A1(_01529_),
    .A2(_01689_),
    .B(_01688_),
    .C(_01690_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08893_ (.I(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08894_ (.A1(_01787_),
    .A2(_01789_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08895_ (.A1(_01784_),
    .A2(_01790_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _08896_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[6] ),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08897_ (.A1(_05280_),
    .A2(_01792_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08898_ (.A1(_06059_),
    .A2(_01791_),
    .B(_01793_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _08899_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[7] ),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08900_ (.A1(_05822_),
    .A2(_01794_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08901_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-19] ),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08902_ (.A1(_01770_),
    .A2(_01773_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08903_ (.A1(_01797_),
    .A2(_01775_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08904_ (.A1(_01709_),
    .A2(_01710_),
    .B(_01708_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08905_ (.A1(_01712_),
    .A2(_01713_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08906_ (.A1(_01799_),
    .A2(_01800_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08907_ (.A1(_01716_),
    .A2(_01767_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08908_ (.A1(_01714_),
    .A2(_01768_),
    .B(_01802_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08909_ (.A1(_01721_),
    .A2(_01735_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08910_ (.A1(_01718_),
    .A2(_01736_),
    .B(_01804_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08911_ (.A1(_06654_),
    .A2(_00373_),
    .A3(_01725_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08912_ (.A1(_01723_),
    .A2(_01724_),
    .B(_01806_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08913_ (.A1(_01805_),
    .A2(_01807_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08914_ (.A1(_06664_),
    .A2(_00370_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08915_ (.A1(_01808_),
    .A2(_01809_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08916_ (.A1(_01740_),
    .A2(_01765_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08917_ (.A1(_01737_),
    .A2(_01766_),
    .B(_01811_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(_01729_),
    .A2(_01733_),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08919_ (.A1(_01726_),
    .A2(_01734_),
    .B(_01813_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08920_ (.A1(_01744_),
    .A2(_01747_),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08921_ (.A1(_01744_),
    .A2(_01747_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08922_ (.A1(_01741_),
    .A2(_01815_),
    .B(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08923_ (.A1(_06659_),
    .A2(_00373_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08924_ (.A1(_06649_),
    .A2(_00379_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08925_ (.A1(_06654_),
    .A2(_00376_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08926_ (.A1(_01819_),
    .A2(_01820_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08927_ (.A1(_01818_),
    .A2(_01821_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08928_ (.A1(_01731_),
    .A2(_01732_),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08929_ (.A1(_01731_),
    .A2(_01732_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08930_ (.A1(_01730_),
    .A2(_01823_),
    .B(_01824_),
    .ZN(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08931_ (.A1(_06642_),
    .A2(_00382_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08932_ (.A1(_06633_),
    .A2(_00388_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08933_ (.A1(_06637_),
    .A2(_00385_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08934_ (.A1(_01826_),
    .A2(_01827_),
    .A3(_01828_),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08935_ (.A1(_01825_),
    .A2(_01829_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08936_ (.A1(_01822_),
    .A2(_01830_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08937_ (.A1(_01814_),
    .A2(_01817_),
    .A3(_01831_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08938_ (.A1(_01750_),
    .A2(_01763_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08939_ (.A1(_01748_),
    .A2(_01764_),
    .B(_01833_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08940_ (.A1(_01745_),
    .A2(_01746_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08941_ (.A1(_01752_),
    .A2(_01753_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08942_ (.A1(_01752_),
    .A2(_01753_),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08943_ (.A1(_01751_),
    .A2(_01836_),
    .B(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08944_ (.A1(_00398_),
    .A2(_06598_),
    .B1(_06618_),
    .B2(_00394_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08945_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06598_),
    .A4(_06618_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08946_ (.A1(_01839_),
    .A2(_01840_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08947_ (.A1(_01835_),
    .A2(_01838_),
    .A3(_01841_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08948_ (.A1(_01757_),
    .A2(_01761_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08949_ (.A1(_01754_),
    .A2(_01762_),
    .B(_01843_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08950_ (.A1(_00355_),
    .A2(_06685_),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08951_ (.A1(_00352_),
    .A2(_06691_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08952_ (.A1(net95),
    .A2(_06627_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08953_ (.A1(_01845_),
    .A2(_01846_),
    .A3(_01847_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08954_ (.A1(net61),
    .A2(_06664_),
    .B1(_06672_),
    .B2(net142),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08955_ (.A1(net61),
    .A2(net142),
    .A3(_06664_),
    .A4(_06672_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08956_ (.A1(_01758_),
    .A2(_01849_),
    .B(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08957_ (.A1(_00357_),
    .A2(_06679_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08958_ (.A1(net158),
    .A2(_06672_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08959_ (.A1(net143),
    .A2(_06674_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08960_ (.A1(_01852_),
    .A2(_01853_),
    .A3(_01854_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08961_ (.A1(_01851_),
    .A2(_01855_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08962_ (.A1(_01848_),
    .A2(_01856_),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08963_ (.A1(_01844_),
    .A2(_01857_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08964_ (.A1(_01842_),
    .A2(_01858_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08965_ (.A1(_01834_),
    .A2(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08966_ (.A1(_01832_),
    .A2(_01860_),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _08967_ (.A1(_01810_),
    .A2(_01812_),
    .A3(_01861_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _08968_ (.A1(_01801_),
    .A2(_01803_),
    .A3(_01862_),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08969_ (.A1(_01706_),
    .A2(_01769_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08970_ (.A1(_01706_),
    .A2(_01769_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08971_ (.A1(_01704_),
    .A2(_01864_),
    .B(_01865_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _08972_ (.A1(_01863_),
    .A2(_01866_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _08973_ (.A1(_01796_),
    .A2(_01798_),
    .A3(_01867_),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08974_ (.A1(_00440_),
    .A2(_01782_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08975_ (.A1(_01869_),
    .A2(_01790_),
    .B(_01783_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08976_ (.A1(_01868_),
    .A2(_01870_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08977_ (.A1(_01868_),
    .A2(_01870_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08978_ (.I(_01872_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08979_ (.A1(_05387_),
    .A2(_01871_),
    .A3(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08980_ (.A1(_01795_),
    .A2(_01874_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08981_ (.I(_01805_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08982_ (.A1(_01875_),
    .A2(_01807_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08983_ (.A1(_06664_),
    .A2(_00370_),
    .A3(_01808_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08984_ (.A1(_01876_),
    .A2(_01877_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08985_ (.A1(_01812_),
    .A2(_01861_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08986_ (.A1(_01812_),
    .A2(_01861_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08987_ (.A1(_01810_),
    .A2(_01879_),
    .B(_01880_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08988_ (.A1(_01817_),
    .A2(_01831_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08989_ (.A1(_01817_),
    .A2(_01831_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08990_ (.A1(_01814_),
    .A2(_01882_),
    .B(_01883_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08991_ (.A1(_06659_),
    .A2(_00373_),
    .A3(_01821_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08992_ (.A1(_01819_),
    .A2(_01820_),
    .B(_01885_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08993_ (.A1(_01884_),
    .A2(_01886_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08994_ (.A1(_00370_),
    .A2(_06672_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08995_ (.A1(_01887_),
    .A2(_01888_),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08996_ (.A1(_01834_),
    .A2(_01859_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08997_ (.A1(_01832_),
    .A2(_01860_),
    .B(_01890_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08998_ (.A1(_01825_),
    .A2(_01829_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08999_ (.A1(_01822_),
    .A2(_01830_),
    .B(_01892_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09000_ (.A1(_01838_),
    .A2(_01841_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09001_ (.A1(_01838_),
    .A2(_01841_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09002_ (.A1(_01835_),
    .A2(_01894_),
    .B(_01895_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09003_ (.A1(_06664_),
    .A2(_00373_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09004_ (.A1(_06654_),
    .A2(_00379_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09005_ (.A1(_06659_),
    .A2(_00376_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09006_ (.A1(_01898_),
    .A2(_01899_),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09007_ (.A1(_01897_),
    .A2(_01900_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09008_ (.A1(_01827_),
    .A2(_01828_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09009_ (.A1(_01827_),
    .A2(_01828_),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09010_ (.A1(_01826_),
    .A2(_01902_),
    .B(_01903_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09011_ (.A1(_06649_),
    .A2(_00382_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09012_ (.A1(_06637_),
    .A2(_00388_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09013_ (.A1(_06642_),
    .A2(_00385_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09014_ (.A1(_01905_),
    .A2(_01906_),
    .A3(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09015_ (.A1(_01904_),
    .A2(_01908_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09016_ (.A1(_01901_),
    .A2(_01909_),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09017_ (.A1(_01893_),
    .A2(_01896_),
    .A3(_01910_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09018_ (.A1(_01844_),
    .A2(_01857_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09019_ (.A1(_01842_),
    .A2(_01858_),
    .B(_01912_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09020_ (.A1(net96),
    .A2(_06627_),
    .B1(_06691_),
    .B2(net138),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09021_ (.A1(net138),
    .A2(net96),
    .A3(_06627_),
    .A4(_06691_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09022_ (.A1(_01845_),
    .A2(_01914_),
    .B(_01915_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09023_ (.A1(_00394_),
    .A2(_06627_),
    .B1(_06618_),
    .B2(_00398_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09024_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06627_),
    .A4(_06618_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09025_ (.A1(_01917_),
    .A2(_01918_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09026_ (.A1(_01916_),
    .A2(_01919_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09027_ (.A1(_01840_),
    .A2(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09028_ (.A1(_01851_),
    .A2(_01855_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09029_ (.A1(_01848_),
    .A2(_01856_),
    .B(_01922_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09030_ (.A1(_00355_),
    .A2(_06691_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09031_ (.A1(net138),
    .A2(_06696_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09032_ (.A1(net95),
    .A2(_06633_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09033_ (.A1(_01924_),
    .A2(_01925_),
    .A3(_01926_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09034_ (.A1(net61),
    .A2(_06672_),
    .B1(_06674_),
    .B2(net60),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09035_ (.A1(net61),
    .A2(net60),
    .A3(_06672_),
    .A4(_06674_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09036_ (.A1(_01852_),
    .A2(_01928_),
    .B(_01929_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09037_ (.A1(_00357_),
    .A2(_06685_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09038_ (.A1(net92),
    .A2(_06674_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09039_ (.A1(net60),
    .A2(_06679_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09040_ (.A1(_01931_),
    .A2(_01932_),
    .A3(_01933_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09041_ (.A1(_01930_),
    .A2(_01934_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09042_ (.A1(_01927_),
    .A2(_01935_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09043_ (.A1(_01921_),
    .A2(_01923_),
    .A3(_01936_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09044_ (.A1(_01937_),
    .A2(_01913_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09045_ (.A1(_01911_),
    .A2(_01938_),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09046_ (.A1(_01891_),
    .A2(_01939_),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09047_ (.A1(_01889_),
    .A2(_01940_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09048_ (.A1(_01881_),
    .A2(_01941_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09049_ (.A1(_01878_),
    .A2(_01942_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09050_ (.A1(_01803_),
    .A2(_01862_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09051_ (.A1(_01803_),
    .A2(_01862_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09052_ (.A1(_01801_),
    .A2(_01944_),
    .B(_01945_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09053_ (.A1(_01943_),
    .A2(_01946_),
    .Z(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09054_ (.A1(_01863_),
    .A2(_01866_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09055_ (.A1(_01797_),
    .A2(_01948_),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09056_ (.A1(_01863_),
    .A2(_01866_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09057_ (.A1(_01775_),
    .A2(_01949_),
    .B(_01950_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09058_ (.A1(_00449_),
    .A2(_01947_),
    .A3(_01951_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09059_ (.A1(_01798_),
    .A2(_01867_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09060_ (.A1(_01796_),
    .A2(_01953_),
    .B(_01873_),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09061_ (.A1(_01952_),
    .A2(_01954_),
    .Z(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _09062_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[8] ),
    .Z(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09063_ (.A1(_05280_),
    .A2(_01956_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09064_ (.A1(_06059_),
    .A2(_01955_),
    .B(_01957_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09065_ (.A1(_01868_),
    .A2(_01952_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _09066_ (.A1(_01788_),
    .A2(_01784_),
    .A3(_01958_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09067_ (.I(_01947_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09068_ (.A1(_01775_),
    .A2(_01949_),
    .B(_01960_),
    .C(_01950_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09069_ (.A1(_01947_),
    .A2(_01951_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09070_ (.A1(_01961_),
    .A2(_01962_),
    .B(_00449_),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09071_ (.A1(_00449_),
    .A2(_01961_),
    .A3(_01962_),
    .B1(_01953_),
    .B2(_01796_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09072_ (.A1(_01787_),
    .A2(_01781_),
    .B(_01868_),
    .C(_01952_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09073_ (.A1(_01963_),
    .A2(_01964_),
    .B1(_01965_),
    .B2(_01783_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09074_ (.A1(_01959_),
    .A2(_01966_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09075_ (.A1(_01943_),
    .A2(_01946_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09076_ (.I(_01968_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09077_ (.A1(_01776_),
    .A2(_01778_),
    .B(_01779_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09078_ (.A1(_01770_),
    .A2(_01773_),
    .B1(_01863_),
    .B2(_01866_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09079_ (.A1(_01863_),
    .A2(_01866_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09080_ (.A1(_01970_),
    .A2(_01971_),
    .B(_01947_),
    .C(_01972_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09081_ (.A1(_01969_),
    .A2(_01973_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09082_ (.A1(_01881_),
    .A2(_01941_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09083_ (.A1(_01878_),
    .A2(_01942_),
    .B(_01975_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09084_ (.I(_01884_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09085_ (.A1(_01977_),
    .A2(_01886_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09086_ (.A1(_01887_),
    .A2(_01888_),
    .B(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09087_ (.A1(_01891_),
    .A2(_01939_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09088_ (.A1(_01889_),
    .A2(_01940_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09089_ (.A1(_01980_),
    .A2(_01981_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09090_ (.A1(_01896_),
    .A2(_01910_),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09091_ (.A1(_01896_),
    .A2(_01910_),
    .Z(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09092_ (.A1(_01893_),
    .A2(_01983_),
    .B(_01984_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09093_ (.A1(_06664_),
    .A2(_00373_),
    .A3(_01900_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09094_ (.A1(_01898_),
    .A2(_01899_),
    .B(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09095_ (.A1(_01985_),
    .A2(_01987_),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09096_ (.A1(_00370_),
    .A2(_06674_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09097_ (.A1(_01988_),
    .A2(_01989_),
    .Z(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09098_ (.A1(_01913_),
    .A2(_01937_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09099_ (.A1(_01911_),
    .A2(net160),
    .B(_01991_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09100_ (.A1(_01904_),
    .A2(_01908_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09101_ (.A1(_01901_),
    .A2(_01909_),
    .B(_01993_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09102_ (.A1(_01916_),
    .A2(_01919_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09103_ (.A1(_01840_),
    .A2(_01920_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09104_ (.A1(_01995_),
    .A2(_01996_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09105_ (.A1(_00373_),
    .A2(_06672_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09106_ (.A1(_06659_),
    .A2(_00379_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09107_ (.A1(_06664_),
    .A2(_00376_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09108_ (.A1(_01999_),
    .A2(_02000_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09109_ (.A1(_01998_),
    .A2(_02001_),
    .Z(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09110_ (.A1(_01906_),
    .A2(_01907_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09111_ (.A1(_01906_),
    .A2(_01907_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09112_ (.A1(_01905_),
    .A2(_02003_),
    .B(_02004_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09113_ (.A1(_06654_),
    .A2(_00382_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09114_ (.A1(_06642_),
    .A2(_00388_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09115_ (.A1(_06649_),
    .A2(_00385_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09116_ (.A1(_02006_),
    .A2(_02007_),
    .A3(_02008_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09117_ (.A1(_02005_),
    .A2(_02009_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09118_ (.A1(_02002_),
    .A2(_02010_),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09119_ (.A1(_01997_),
    .A2(_02011_),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09120_ (.A1(_01994_),
    .A2(_02012_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09121_ (.A1(_01923_),
    .A2(_01936_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09122_ (.A1(_01923_),
    .A2(_01936_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09123_ (.A1(_01921_),
    .A2(_02014_),
    .B(_02015_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09124_ (.A1(net96),
    .A2(_06633_),
    .B1(_06696_),
    .B2(net137),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09125_ (.A1(net137),
    .A2(net96),
    .A3(_06633_),
    .A4(_06696_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09126_ (.A1(_01924_),
    .A2(_02017_),
    .B(_02018_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09127_ (.A1(_00398_),
    .A2(_06627_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09128_ (.A1(_06633_),
    .A2(_00394_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09129_ (.A1(_02020_),
    .A2(_02021_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09130_ (.A1(_02019_),
    .A2(_02022_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09131_ (.A1(_01918_),
    .A2(_02023_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09132_ (.A1(_01930_),
    .A2(_01934_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09133_ (.A1(_01927_),
    .A2(_01935_),
    .B(_02025_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09134_ (.A1(_00355_),
    .A2(_06696_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09135_ (.A1(net58),
    .A2(_06701_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09136_ (.A1(_06637_),
    .A2(net95),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09137_ (.A1(_02027_),
    .A2(_02028_),
    .A3(_02029_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09138_ (.A1(net61),
    .A2(_06674_),
    .B1(_06679_),
    .B2(net60),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09139_ (.A1(net61),
    .A2(net60),
    .A3(_06674_),
    .A4(_06679_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09140_ (.A1(_01931_),
    .A2(_02031_),
    .B(_02032_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09141_ (.A1(net73),
    .A2(_06691_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09142_ (.A1(net61),
    .A2(_06679_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09143_ (.A1(net60),
    .A2(_06685_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09144_ (.A1(_02034_),
    .A2(_02035_),
    .A3(_02036_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09145_ (.A1(_02033_),
    .A2(_02037_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09146_ (.A1(_02030_),
    .A2(_02038_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09147_ (.A1(_02024_),
    .A2(_02026_),
    .A3(_02039_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09148_ (.A1(_02016_),
    .A2(_02040_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09149_ (.A1(_02013_),
    .A2(_02041_),
    .Z(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09150_ (.A1(_01992_),
    .A2(_02042_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09151_ (.A1(_01990_),
    .A2(_02043_),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09152_ (.I(_02044_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09153_ (.A1(_01979_),
    .A2(_01982_),
    .A3(_02045_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09154_ (.A1(_02046_),
    .A2(_01976_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09155_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-17] ),
    .A2(_01974_),
    .A3(_02047_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09156_ (.A1(_01967_),
    .A2(_02048_),
    .Z(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09157_ (.A1(_01967_),
    .A2(_02048_),
    .B(_05182_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _09158_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[9] ),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09159_ (.A1(_05280_),
    .A2(_02051_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09160_ (.A1(_02049_),
    .A2(_02050_),
    .B(_02052_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09161_ (.A1(_01774_),
    .A2(_01867_),
    .A3(_01947_),
    .A4(_02047_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09162_ (.A1(_01700_),
    .A2(_02053_),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09163_ (.A1(_01513_),
    .A2(_01518_),
    .B(_02054_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09164_ (.I(_02046_),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09165_ (.A1(_01976_),
    .A2(_02056_),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09166_ (.A1(_01972_),
    .A2(_01947_),
    .A3(_01971_),
    .A4(_02047_),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09167_ (.A1(_01976_),
    .A2(_02056_),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09168_ (.A1(_01969_),
    .A2(_02057_),
    .B(_02058_),
    .C(_02059_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09169_ (.A1(_01695_),
    .A2(_01698_),
    .B(_02053_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09170_ (.A1(_02060_),
    .A2(_02061_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09171_ (.I(_01985_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09172_ (.A1(_02063_),
    .A2(_01987_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09173_ (.A1(_01988_),
    .A2(_01989_),
    .B(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09174_ (.A1(_01992_),
    .A2(_02042_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09175_ (.A1(_01990_),
    .A2(_02043_),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09176_ (.A1(_02066_),
    .A2(_02067_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09177_ (.A1(_01997_),
    .A2(_02011_),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09178_ (.A1(_01994_),
    .A2(_02012_),
    .B(_02069_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09179_ (.A1(_00373_),
    .A2(_06672_),
    .A3(_02001_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09180_ (.A1(_01999_),
    .A2(_02000_),
    .B(_02071_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09181_ (.A1(_02070_),
    .A2(_02072_),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09182_ (.A1(_00370_),
    .A2(_06679_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09183_ (.A1(_02073_),
    .A2(_02074_),
    .Z(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09184_ (.A1(_02016_),
    .A2(_02040_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09185_ (.A1(_02013_),
    .A2(_02041_),
    .B(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09186_ (.A1(_02005_),
    .A2(_02009_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09187_ (.A1(_02002_),
    .A2(_02010_),
    .B(_02078_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09188_ (.A1(_02019_),
    .A2(_02022_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09189_ (.A1(_01918_),
    .A2(_02023_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09190_ (.A1(_02080_),
    .A2(_02081_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09191_ (.A1(_00373_),
    .A2(_06674_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09192_ (.A1(_06664_),
    .A2(_00379_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09193_ (.A1(_00376_),
    .A2(_06672_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09194_ (.A1(_02084_),
    .A2(_02085_),
    .Z(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09195_ (.A1(_02083_),
    .A2(_02086_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09196_ (.A1(_02007_),
    .A2(_02008_),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09197_ (.A1(_02007_),
    .A2(_02008_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09198_ (.A1(_02006_),
    .A2(_02088_),
    .B(_02089_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09199_ (.A1(_06659_),
    .A2(_00382_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09200_ (.A1(_06649_),
    .A2(_00388_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09201_ (.A1(_06654_),
    .A2(_00385_),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09202_ (.A1(_02091_),
    .A2(_02092_),
    .A3(_02093_),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09203_ (.A1(_02090_),
    .A2(_02094_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09204_ (.A1(_02087_),
    .A2(_02095_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09205_ (.A1(_02082_),
    .A2(_02096_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09206_ (.A1(_02079_),
    .A2(_02097_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09207_ (.A1(_02026_),
    .A2(_02039_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09208_ (.A1(_02026_),
    .A2(_02039_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09209_ (.A1(_02024_),
    .A2(_02099_),
    .B(_02100_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09210_ (.A1(_02020_),
    .A2(_02021_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09211_ (.A1(_02028_),
    .A2(_02029_),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09212_ (.A1(_02028_),
    .A2(_02029_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09213_ (.A1(_02027_),
    .A2(_02103_),
    .B(_02104_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09214_ (.A1(_06633_),
    .A2(_00398_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09215_ (.A1(_06637_),
    .A2(_00394_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09216_ (.A1(_02106_),
    .A2(_02107_),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09217_ (.A1(_02102_),
    .A2(_02105_),
    .A3(_02108_),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09218_ (.A1(_02033_),
    .A2(_02037_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09219_ (.A1(_02030_),
    .A2(_02038_),
    .B(_02110_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09220_ (.A1(_00355_),
    .A2(_06701_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09221_ (.A1(_06642_),
    .A2(net98),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09222_ (.A1(net58),
    .A2(_06708_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09223_ (.A1(_02112_),
    .A2(_02113_),
    .A3(_02114_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09224_ (.A1(net61),
    .A2(_06679_),
    .B1(_06685_),
    .B2(net60),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09225_ (.A1(net61),
    .A2(net60),
    .A3(_06679_),
    .A4(_06685_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09226_ (.A1(_02034_),
    .A2(_02116_),
    .B(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09227_ (.A1(net73),
    .A2(_06696_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09228_ (.A1(net91),
    .A2(_06685_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09229_ (.A1(net60),
    .A2(_06691_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09230_ (.A1(_02119_),
    .A2(_02120_),
    .A3(_02121_),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09231_ (.A1(_02118_),
    .A2(_02122_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09232_ (.A1(_02115_),
    .A2(_02123_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09233_ (.A1(_02111_),
    .A2(_02124_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09234_ (.A1(_02109_),
    .A2(_02125_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09235_ (.A1(_02101_),
    .A2(_02126_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09236_ (.A1(_02098_),
    .A2(_02127_),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09237_ (.A1(_02077_),
    .A2(_02128_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09238_ (.A1(_02075_),
    .A2(_02129_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09239_ (.I(_02130_),
    .ZN(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09240_ (.A1(_02068_),
    .A2(_02131_),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09241_ (.A1(_02065_),
    .A2(_02132_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09242_ (.A1(_01982_),
    .A2(_02045_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09243_ (.A1(_01980_),
    .A2(_01981_),
    .A3(_02044_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09244_ (.A1(_01979_),
    .A2(_02134_),
    .A3(_02135_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09245_ (.A1(_02134_),
    .A2(_02136_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09246_ (.A1(_02133_),
    .A2(_02137_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09247_ (.A1(_02055_),
    .A2(_02062_),
    .B(_02138_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09248_ (.I(_02138_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09249_ (.A1(net56),
    .A2(_01348_),
    .B(_01700_),
    .C(_02053_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09250_ (.A1(_02060_),
    .A2(_02061_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09251_ (.A1(_02140_),
    .A2(_02141_),
    .A3(_02142_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09252_ (.A1(_02139_),
    .A2(_02143_),
    .Z(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09253_ (.A1(_00459_),
    .A2(_02144_),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09254_ (.A1(_01976_),
    .A2(_02056_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09255_ (.A1(_01968_),
    .A2(_01961_),
    .B1(_02146_),
    .B2(_02057_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09256_ (.A1(_01969_),
    .A2(_01973_),
    .A3(_02047_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09257_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-17] ),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09258_ (.A1(_02147_),
    .A2(_02148_),
    .B(_02149_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09259_ (.A1(_02150_),
    .A2(_02049_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09260_ (.A1(_02145_),
    .A2(_02151_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _09261_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[10] ),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09262_ (.A1(_05280_),
    .A2(_02153_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09263_ (.A1(_06059_),
    .A2(_02152_),
    .B(_02154_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09264_ (.A1(_02134_),
    .A2(_02136_),
    .B(_02133_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09265_ (.A1(_02155_),
    .A2(_02139_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09266_ (.A1(_02068_),
    .A2(_02131_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09267_ (.A1(_02065_),
    .A2(_02132_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09268_ (.I(_02070_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09269_ (.A1(_02159_),
    .A2(_02072_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09270_ (.A1(_02073_),
    .A2(_02074_),
    .B(_02160_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09271_ (.A1(_02077_),
    .A2(_02128_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09272_ (.A1(_02075_),
    .A2(_02129_),
    .B(_02162_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09273_ (.A1(_02082_),
    .A2(_02096_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09274_ (.A1(_02079_),
    .A2(_02097_),
    .B(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09275_ (.A1(_00373_),
    .A2(_06674_),
    .A3(_02086_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09276_ (.A1(_02084_),
    .A2(_02085_),
    .B(_02166_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09277_ (.A1(_02165_),
    .A2(_02167_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09278_ (.A1(_00370_),
    .A2(_06685_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09279_ (.A1(_02168_),
    .A2(_02169_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09280_ (.A1(_02101_),
    .A2(_02126_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09281_ (.A1(_02098_),
    .A2(_02127_),
    .B(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09282_ (.A1(_02090_),
    .A2(_02094_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09283_ (.A1(_02087_),
    .A2(_02095_),
    .B(_02173_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09284_ (.A1(_02105_),
    .A2(_02108_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09285_ (.A1(_02105_),
    .A2(_02108_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09286_ (.A1(_02102_),
    .A2(_02175_),
    .B(_02176_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09287_ (.A1(_00373_),
    .A2(_06679_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09288_ (.A1(_00379_),
    .A2(_06672_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09289_ (.A1(_00376_),
    .A2(_06674_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09290_ (.A1(_02179_),
    .A2(_02180_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09291_ (.A1(_02178_),
    .A2(_02181_),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09292_ (.A1(_02092_),
    .A2(_02093_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09293_ (.A1(_02092_),
    .A2(_02093_),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09294_ (.A1(_02091_),
    .A2(_02183_),
    .B(_02184_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09295_ (.A1(_06664_),
    .A2(_00382_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09296_ (.A1(_06654_),
    .A2(_00388_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09297_ (.A1(_06659_),
    .A2(_00385_),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09298_ (.A1(_02186_),
    .A2(_02187_),
    .A3(_02188_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09299_ (.A1(_02185_),
    .A2(_02189_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09300_ (.A1(_02182_),
    .A2(_02190_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09301_ (.A1(_02174_),
    .A2(_02177_),
    .A3(_02191_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09302_ (.A1(_02111_),
    .A2(_02124_),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09303_ (.A1(_02109_),
    .A2(_02125_),
    .B(_02193_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09304_ (.A1(_02106_),
    .A2(_02107_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09305_ (.A1(_02113_),
    .A2(_02114_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09306_ (.A1(_02113_),
    .A2(_02114_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09307_ (.A1(_02112_),
    .A2(_02196_),
    .B(_02197_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09308_ (.A1(_06637_),
    .A2(_00398_),
    .B1(_00394_),
    .B2(_06642_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09309_ (.A1(_06642_),
    .A2(_06637_),
    .A3(_00398_),
    .A4(_00394_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09310_ (.A1(_02199_),
    .A2(_02200_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09311_ (.A1(_02195_),
    .A2(_02198_),
    .A3(_02201_),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09312_ (.A1(_02118_),
    .A2(_02122_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09313_ (.A1(_02115_),
    .A2(_02123_),
    .B(_02203_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09314_ (.A1(net61),
    .A2(_06685_),
    .B1(_06691_),
    .B2(net60),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09315_ (.A1(net61),
    .A2(net60),
    .A3(_06685_),
    .A4(_06691_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09316_ (.A1(_02119_),
    .A2(_02205_),
    .B(_02206_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09317_ (.A1(_00357_),
    .A2(_06701_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09318_ (.A1(net91),
    .A2(_06691_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09319_ (.A1(net60),
    .A2(_06696_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09320_ (.A1(_02208_),
    .A2(_02209_),
    .A3(_02210_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09321_ (.A1(_02207_),
    .A2(_02211_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09322_ (.A1(_00355_),
    .A2(_06708_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09323_ (.A1(net137),
    .A2(_06710_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09324_ (.A1(_06649_),
    .A2(net95),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09325_ (.A1(_02213_),
    .A2(_02214_),
    .A3(_02215_),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09326_ (.A1(_02212_),
    .A2(_02216_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09327_ (.A1(_02204_),
    .A2(_02217_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09328_ (.A1(_02202_),
    .A2(_02218_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09329_ (.A1(_02194_),
    .A2(_02219_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09330_ (.A1(_02192_),
    .A2(_02220_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09331_ (.A1(_02172_),
    .A2(_02221_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09332_ (.A1(_02170_),
    .A2(_02222_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _09333_ (.A1(_02161_),
    .A2(_02163_),
    .A3(_02223_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09334_ (.A1(_02157_),
    .A2(_02158_),
    .B(_02224_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09335_ (.A1(_02157_),
    .A2(_02158_),
    .A3(_02224_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09336_ (.A1(_02225_),
    .A2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09337_ (.A1(_02156_),
    .A2(_02227_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09338_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-15] ),
    .A2(_02228_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09339_ (.A1(_00459_),
    .A2(_02144_),
    .ZN(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09340_ (.A1(_00459_),
    .A2(_02144_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09341_ (.A1(_02150_),
    .A2(_02049_),
    .A3(_02230_),
    .B(_02231_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09342_ (.A1(_02229_),
    .A2(_02232_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09343_ (.A1(_02229_),
    .A2(_02232_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09344_ (.A1(_05182_),
    .A2(_02234_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _09345_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[11] ),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09346_ (.A1(_05280_),
    .A2(_02236_),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09347_ (.A1(_02233_),
    .A2(_02235_),
    .B(_02237_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _09348_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[12] ),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09349_ (.I(_02165_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09350_ (.A1(_02239_),
    .A2(_02167_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09351_ (.A1(_02168_),
    .A2(_02169_),
    .B(_02240_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09352_ (.A1(_02172_),
    .A2(_02221_),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09353_ (.A1(_02170_),
    .A2(_02222_),
    .B(_02242_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09354_ (.A1(_02177_),
    .A2(_02191_),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09355_ (.A1(_02177_),
    .A2(_02191_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09356_ (.A1(_02174_),
    .A2(_02244_),
    .B(_02245_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09357_ (.A1(_00373_),
    .A2(_06679_),
    .A3(_02181_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09358_ (.A1(_02179_),
    .A2(_02180_),
    .B(_02247_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09359_ (.A1(_02246_),
    .A2(_02248_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09360_ (.A1(_00370_),
    .A2(_06691_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09361_ (.A1(_02249_),
    .A2(_02250_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09362_ (.A1(_02194_),
    .A2(_02219_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09363_ (.A1(_02192_),
    .A2(_02220_),
    .B(_02252_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09364_ (.A1(_02185_),
    .A2(_02189_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09365_ (.A1(_02182_),
    .A2(_02190_),
    .B(_02254_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09366_ (.A1(_02198_),
    .A2(_02201_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09367_ (.A1(_02198_),
    .A2(_02201_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09368_ (.A1(_02195_),
    .A2(_02256_),
    .B(_02257_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09369_ (.A1(_00373_),
    .A2(_06685_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09370_ (.A1(_00379_),
    .A2(_06674_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09371_ (.A1(_00376_),
    .A2(_06679_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09372_ (.A1(_02260_),
    .A2(_02261_),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09373_ (.A1(_02259_),
    .A2(_02262_),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09374_ (.A1(_02187_),
    .A2(_02188_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09375_ (.A1(_02187_),
    .A2(_02188_),
    .Z(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09376_ (.A1(_02186_),
    .A2(_02264_),
    .B(_02265_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09377_ (.A1(_00382_),
    .A2(_06672_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09378_ (.A1(_06659_),
    .A2(_00388_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09379_ (.A1(_06664_),
    .A2(_00385_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09380_ (.A1(_02267_),
    .A2(_02268_),
    .A3(_02269_),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09381_ (.A1(_02266_),
    .A2(_02270_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09382_ (.A1(_02263_),
    .A2(_02271_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09383_ (.A1(_02255_),
    .A2(_02258_),
    .A3(_02272_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09384_ (.A1(_02204_),
    .A2(_02217_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09385_ (.A1(_02202_),
    .A2(_02218_),
    .B(_02274_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09386_ (.A1(_02207_),
    .A2(_02211_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09387_ (.A1(_02212_),
    .A2(_02216_),
    .B(_02276_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09388_ (.A1(net61),
    .A2(_06691_),
    .B1(_06696_),
    .B2(net142),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09389_ (.A1(net61),
    .A2(net142),
    .A3(_06691_),
    .A4(_06696_),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09390_ (.A1(_02208_),
    .A2(_02278_),
    .B(_02279_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09391_ (.A1(_00357_),
    .A2(_06708_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09392_ (.A1(net92),
    .A2(_06696_),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09393_ (.A1(net142),
    .A2(_06701_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09394_ (.A1(_02281_),
    .A2(_02282_),
    .A3(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09395_ (.A1(_02280_),
    .A2(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09396_ (.A1(_00355_),
    .A2(_06710_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09397_ (.A1(_06654_),
    .A2(net96),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09398_ (.A1(net58),
    .A2(_06724_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09399_ (.A1(_02286_),
    .A2(_02287_),
    .A3(_02288_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09400_ (.A1(_02285_),
    .A2(_02289_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09401_ (.A1(_02277_),
    .A2(_02290_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09402_ (.A1(_06649_),
    .A2(net95),
    .B1(_06710_),
    .B2(net58),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09403_ (.A1(_06649_),
    .A2(net58),
    .A3(net95),
    .A4(_06710_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09404_ (.A1(_02213_),
    .A2(_02292_),
    .B(_02293_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09405_ (.A1(_06642_),
    .A2(_00398_),
    .B1(_00394_),
    .B2(_06649_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09406_ (.A1(_06642_),
    .A2(_06649_),
    .A3(_00398_),
    .A4(_00394_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09407_ (.A1(_02295_),
    .A2(_02296_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09408_ (.A1(_02294_),
    .A2(_02297_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09409_ (.A1(_02200_),
    .A2(_02298_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09410_ (.A1(_02291_),
    .A2(_02299_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09411_ (.A1(_02275_),
    .A2(_02300_),
    .Z(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09412_ (.A1(_02273_),
    .A2(_02301_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09413_ (.A1(_02253_),
    .A2(_02302_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09414_ (.A1(_02251_),
    .A2(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09415_ (.A1(_02243_),
    .A2(_02304_),
    .Z(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09416_ (.A1(_02241_),
    .A2(_02305_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09417_ (.A1(_02163_),
    .A2(_02223_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09418_ (.A1(_02163_),
    .A2(_02223_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09419_ (.A1(_02161_),
    .A2(_02307_),
    .B(_02308_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09420_ (.A1(_02306_),
    .A2(_02309_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09421_ (.A1(_02157_),
    .A2(_02158_),
    .A3(_02224_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _09422_ (.A1(_02155_),
    .A2(_02139_),
    .A3(_02225_),
    .B(_02311_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09423_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-14] ),
    .A2(_02310_),
    .A3(_02312_),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09424_ (.A1(_00463_),
    .A2(_02228_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09425_ (.A1(_02314_),
    .A2(_02233_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09426_ (.A1(_02313_),
    .A2(_02315_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09427_ (.I0(_02238_),
    .I1(_02316_),
    .S(_00395_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09428_ (.I(_02317_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09429_ (.A1(_02306_),
    .A2(_02309_),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09430_ (.A1(_02310_),
    .A2(_02312_),
    .B(_02318_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09431_ (.A1(_02243_),
    .A2(_02304_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09432_ (.A1(_02241_),
    .A2(_02305_),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09433_ (.I(_02246_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09434_ (.A1(_02322_),
    .A2(_02248_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09435_ (.A1(_00370_),
    .A2(_06691_),
    .A3(_02249_),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09436_ (.A1(_02323_),
    .A2(_02324_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09437_ (.A1(_02253_),
    .A2(_02302_),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09438_ (.A1(_02251_),
    .A2(_02303_),
    .B(_02326_),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09439_ (.A1(_02258_),
    .A2(_02272_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09440_ (.A1(_02258_),
    .A2(_02272_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09441_ (.A1(_02255_),
    .A2(_02328_),
    .B(_02329_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09442_ (.A1(_00373_),
    .A2(_06685_),
    .A3(_02262_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09443_ (.A1(_02260_),
    .A2(_02261_),
    .B(_02331_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09444_ (.A1(_02330_),
    .A2(_02332_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09445_ (.A1(_00370_),
    .A2(_06696_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09446_ (.A1(_02333_),
    .A2(_02334_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09447_ (.A1(_02202_),
    .A2(_02218_),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09448_ (.A1(_02274_),
    .A2(_02336_),
    .B(_02300_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09449_ (.A1(_02273_),
    .A2(_02301_),
    .B(_02337_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09450_ (.A1(_02277_),
    .A2(_02290_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09451_ (.A1(_02291_),
    .A2(_02299_),
    .B(_02339_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09452_ (.A1(_02280_),
    .A2(_02284_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09453_ (.A1(_02285_),
    .A2(_02289_),
    .B(_02341_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09454_ (.A1(net91),
    .A2(_06696_),
    .B1(_06701_),
    .B2(net142),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09455_ (.A1(net91),
    .A2(net142),
    .A3(_06696_),
    .A4(_06701_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09456_ (.A1(_02281_),
    .A2(_02343_),
    .B(_02344_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09457_ (.A1(_00357_),
    .A2(_06710_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09458_ (.A1(net158),
    .A2(_06701_),
    .ZN(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09459_ (.A1(net142),
    .A2(_06708_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09460_ (.A1(_02346_),
    .A2(_02347_),
    .A3(_02348_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09461_ (.A1(_02345_),
    .A2(_02349_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09462_ (.A1(_00355_),
    .A2(_06724_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09463_ (.A1(net96),
    .A2(_06659_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09464_ (.A1(net137),
    .A2(_06730_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09465_ (.A1(_02351_),
    .A2(_02352_),
    .A3(_02353_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09466_ (.A1(_02350_),
    .A2(_02354_),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09467_ (.A1(_02342_),
    .A2(_02355_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09468_ (.A1(_06654_),
    .A2(net95),
    .B1(_06724_),
    .B2(net58),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09469_ (.A1(_06654_),
    .A2(net58),
    .A3(net95),
    .A4(_06724_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09470_ (.A1(_02286_),
    .A2(_02357_),
    .B(_02358_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09471_ (.A1(_06649_),
    .A2(_00398_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09472_ (.A1(_06654_),
    .A2(_00394_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09473_ (.A1(_02360_),
    .A2(_02361_),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09474_ (.A1(_02359_),
    .A2(_02362_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09475_ (.A1(_02296_),
    .A2(_02363_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09476_ (.A1(_02340_),
    .A2(_02356_),
    .A3(_02364_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09477_ (.A1(_02266_),
    .A2(_02270_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09478_ (.A1(_02263_),
    .A2(_02271_),
    .B(_02366_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09479_ (.A1(_02294_),
    .A2(_02297_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09480_ (.A1(_02200_),
    .A2(_02298_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09481_ (.A1(_02368_),
    .A2(_02369_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09482_ (.A1(_00373_),
    .A2(_06691_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09483_ (.A1(_00379_),
    .A2(_06679_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09484_ (.A1(_00376_),
    .A2(_06685_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09485_ (.A1(_02372_),
    .A2(_02373_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09486_ (.A1(_02371_),
    .A2(_02374_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09487_ (.A1(_02268_),
    .A2(_02269_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09488_ (.A1(_02268_),
    .A2(_02269_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09489_ (.A1(_02267_),
    .A2(_02376_),
    .B(_02377_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(_00382_),
    .A2(_06674_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09491_ (.A1(_06664_),
    .A2(_00388_),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09492_ (.A1(_00385_),
    .A2(_06672_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09493_ (.A1(_02379_),
    .A2(_02380_),
    .A3(_02381_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09494_ (.A1(_02378_),
    .A2(_02382_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09495_ (.A1(_02375_),
    .A2(_02383_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09496_ (.A1(_02370_),
    .A2(_02384_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09497_ (.A1(_02367_),
    .A2(_02385_),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09498_ (.A1(_02365_),
    .A2(_02386_),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09499_ (.A1(_02338_),
    .A2(_02387_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09500_ (.A1(_02335_),
    .A2(_02388_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09501_ (.A1(_02325_),
    .A2(_02327_),
    .A3(_02389_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09502_ (.A1(_02320_),
    .A2(_02321_),
    .B(_02390_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _09503_ (.A1(_02320_),
    .A2(_02321_),
    .A3(_02390_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09504_ (.A1(_02391_),
    .A2(_02392_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09505_ (.A1(_02319_),
    .A2(_02393_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09506_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-13] ),
    .A2(_02394_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09507_ (.A1(_00463_),
    .A2(_02156_),
    .A3(_02227_),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09508_ (.A1(_02396_),
    .A2(_02313_),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09509_ (.A1(_02048_),
    .A2(_02145_),
    .A3(_02397_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09510_ (.A1(_02150_),
    .A2(_02230_),
    .B(_02231_),
    .C(_02397_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09511_ (.A1(_02310_),
    .A2(_02312_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09512_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-14] ),
    .A2(_02400_),
    .Z(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09513_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-14] ),
    .A2(_02400_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09514_ (.A1(_02314_),
    .A2(_02401_),
    .B(_02402_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09515_ (.A1(_02399_),
    .A2(_02403_),
    .ZN(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09516_ (.A1(_01967_),
    .A2(_02398_),
    .B(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09517_ (.A1(_02395_),
    .A2(_02405_),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09518_ (.A1(_02395_),
    .A2(_02405_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09519_ (.A1(_05182_),
    .A2(_02407_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _09520_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[13] ),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09521_ (.A1(_05280_),
    .A2(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09522_ (.A1(_02406_),
    .A2(_02408_),
    .B(_02410_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09523_ (.I(_02330_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09524_ (.A1(_02411_),
    .A2(_02332_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09525_ (.A1(_00370_),
    .A2(_06696_),
    .A3(_02333_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09526_ (.A1(_02412_),
    .A2(_02413_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09527_ (.A1(_02338_),
    .A2(_02387_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09528_ (.A1(_02335_),
    .A2(_02388_),
    .B(_02415_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09529_ (.A1(_02356_),
    .A2(_02364_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09530_ (.A1(_02356_),
    .A2(_02364_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09531_ (.A1(_02340_),
    .A2(_02417_),
    .A3(_02418_),
    .B1(_02365_),
    .B2(_02386_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09532_ (.A1(_02342_),
    .A2(_02355_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09533_ (.A1(_02356_),
    .A2(_02364_),
    .B(_02420_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09534_ (.A1(_02345_),
    .A2(_02349_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09535_ (.A1(_02350_),
    .A2(_02354_),
    .B(_02422_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09536_ (.A1(net61),
    .A2(_06701_),
    .B1(_06708_),
    .B2(net142),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09537_ (.A1(net61),
    .A2(net142),
    .A3(_06701_),
    .A4(_06708_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09538_ (.A1(_02346_),
    .A2(_02424_),
    .B(_02425_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09539_ (.A1(_00357_),
    .A2(_06724_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09540_ (.A1(net92),
    .A2(_06708_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09541_ (.A1(net142),
    .A2(_06710_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09542_ (.A1(_02427_),
    .A2(_02428_),
    .A3(_02429_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09543_ (.A1(_02426_),
    .A2(_02430_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09544_ (.A1(_00355_),
    .A2(_06730_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09545_ (.A1(_06664_),
    .A2(net96),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09546_ (.A1(net137),
    .A2(_06738_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09547_ (.A1(_02432_),
    .A2(_02433_),
    .A3(_02434_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09548_ (.A1(_02431_),
    .A2(_02435_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09549_ (.A1(_02423_),
    .A2(_02436_),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09550_ (.A1(_02360_),
    .A2(_02361_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09551_ (.A1(_02352_),
    .A2(_02353_),
    .Z(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09552_ (.A1(_02352_),
    .A2(_02353_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09553_ (.A1(_02351_),
    .A2(_02439_),
    .B(_02440_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09554_ (.A1(_06654_),
    .A2(_00398_),
    .B1(_00394_),
    .B2(_06659_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09555_ (.A1(_06654_),
    .A2(_06659_),
    .A3(_00398_),
    .A4(_00394_),
    .Z(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09556_ (.A1(_02442_),
    .A2(_02443_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09557_ (.A1(_02438_),
    .A2(_02441_),
    .A3(_02444_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09558_ (.A1(_02421_),
    .A2(_02437_),
    .A3(_02445_),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09559_ (.A1(_02378_),
    .A2(_02382_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09560_ (.A1(_02375_),
    .A2(_02383_),
    .B(_02447_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09561_ (.A1(_02359_),
    .A2(_02362_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09562_ (.A1(_02296_),
    .A2(_02363_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09563_ (.A1(_02449_),
    .A2(_02450_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09564_ (.A1(_00373_),
    .A2(_06696_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09565_ (.A1(_00379_),
    .A2(_06685_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09566_ (.A1(_00376_),
    .A2(_06691_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09567_ (.A1(_02453_),
    .A2(_02454_),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09568_ (.A1(_02452_),
    .A2(_02455_),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09569_ (.A1(_02380_),
    .A2(_02381_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09570_ (.A1(_02380_),
    .A2(_02381_),
    .Z(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09571_ (.A1(_02379_),
    .A2(_02457_),
    .B(_02458_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09572_ (.A1(_00382_),
    .A2(_06679_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09573_ (.A1(_00388_),
    .A2(_06672_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09574_ (.A1(_00385_),
    .A2(_06674_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09575_ (.A1(_02460_),
    .A2(_02461_),
    .A3(_02462_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09576_ (.A1(_02459_),
    .A2(_02463_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09577_ (.A1(_02456_),
    .A2(_02464_),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09578_ (.A1(_02451_),
    .A2(_02465_),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09579_ (.A1(_02448_),
    .A2(_02466_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09580_ (.A1(_02446_),
    .A2(_02467_),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09581_ (.A1(_02419_),
    .A2(_02468_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09582_ (.A1(_02370_),
    .A2(_02384_),
    .Z(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09583_ (.A1(_02367_),
    .A2(_02385_),
    .B(_02470_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09584_ (.A1(_00373_),
    .A2(_06691_),
    .A3(_02374_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09585_ (.A1(_02372_),
    .A2(_02373_),
    .B(_02472_),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09586_ (.A1(_02471_),
    .A2(_02473_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09587_ (.A1(_00370_),
    .A2(_06701_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09588_ (.A1(_02474_),
    .A2(_02475_),
    .Z(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09589_ (.A1(_02469_),
    .A2(_02476_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09590_ (.A1(_02416_),
    .A2(_02477_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09591_ (.A1(_02414_),
    .A2(_02478_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09592_ (.I(_02327_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09593_ (.A1(_02480_),
    .A2(_02389_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09594_ (.A1(_02480_),
    .A2(_02389_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09595_ (.A1(_02325_),
    .A2(_02481_),
    .B(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09596_ (.A1(_02479_),
    .A2(_02483_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09597_ (.A1(_02479_),
    .A2(_02483_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09598_ (.A1(_02484_),
    .A2(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09599_ (.I(_02310_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09600_ (.A1(_02227_),
    .A2(_02487_),
    .A3(_02393_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09601_ (.A1(_02055_),
    .A2(_02062_),
    .B(_02488_),
    .C(_02138_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09602_ (.A1(_02487_),
    .A2(_02393_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09603_ (.A1(_02155_),
    .A2(_02225_),
    .B(_02311_),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09604_ (.I(_02391_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09605_ (.A1(_02318_),
    .A2(_02392_),
    .B1(_02490_),
    .B2(_02491_),
    .C(_02492_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09606_ (.A1(_02489_),
    .A2(_02493_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09607_ (.A1(_02486_),
    .A2(_02494_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09608_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-12] ),
    .A2(_02495_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09609_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-13] ),
    .A2(_02394_),
    .B(_02406_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09610_ (.A1(_02496_),
    .A2(_02497_),
    .Z(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _09611_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[14] ),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09612_ (.A1(_05280_),
    .A2(_02499_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09613_ (.A1(_06059_),
    .A2(_02498_),
    .B(_02500_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09614_ (.A1(_02486_),
    .A2(_02494_),
    .B(_02484_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09615_ (.A1(_02416_),
    .A2(_02477_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09616_ (.A1(_02414_),
    .A2(_02478_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09617_ (.I(_02471_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09618_ (.A1(_02504_),
    .A2(_02473_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09619_ (.A1(_02474_),
    .A2(_02475_),
    .B(_02505_),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09620_ (.A1(_02419_),
    .A2(_02468_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09621_ (.A1(_02469_),
    .A2(_02476_),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09622_ (.A1(_02507_),
    .A2(_02508_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09623_ (.A1(_02437_),
    .A2(_02445_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09624_ (.A1(_02437_),
    .A2(_02445_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09625_ (.A1(_02421_),
    .A2(_02510_),
    .A3(_02511_),
    .B1(_02446_),
    .B2(_02467_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09626_ (.A1(_02423_),
    .A2(_02436_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09627_ (.A1(_02437_),
    .A2(_02445_),
    .B(_02513_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09628_ (.A1(_02426_),
    .A2(_02430_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09629_ (.A1(_02431_),
    .A2(_02435_),
    .B(_02515_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09630_ (.A1(net91),
    .A2(_06708_),
    .B1(_06710_),
    .B2(net142),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09631_ (.A1(net91),
    .A2(net142),
    .A3(_06708_),
    .A4(_06710_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09632_ (.A1(_02427_),
    .A2(_02517_),
    .B(_02518_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09633_ (.A1(_00357_),
    .A2(_06730_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09634_ (.A1(net158),
    .A2(_06710_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09635_ (.A1(net143),
    .A2(_06724_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09636_ (.A1(_02520_),
    .A2(_02521_),
    .A3(_02522_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09637_ (.A1(_02519_),
    .A2(_02523_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09638_ (.A1(_00355_),
    .A2(_06738_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09639_ (.A1(net96),
    .A2(_06672_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09640_ (.A1(net138),
    .A2(_06742_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09641_ (.A1(_02525_),
    .A2(_02526_),
    .A3(_02527_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09642_ (.A1(_02524_),
    .A2(_02528_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09643_ (.A1(_02516_),
    .A2(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09644_ (.A1(_02433_),
    .A2(_02434_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09645_ (.A1(_02433_),
    .A2(_02434_),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09646_ (.A1(_02432_),
    .A2(_02531_),
    .B(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09647_ (.A1(_06659_),
    .A2(_00398_),
    .B1(_00394_),
    .B2(_06664_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09648_ (.A1(_06664_),
    .A2(_06659_),
    .A3(_00398_),
    .A4(_00394_),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09649_ (.A1(_02534_),
    .A2(_02535_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09650_ (.A1(_02533_),
    .A2(_02536_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09651_ (.A1(_02443_),
    .A2(_02537_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09652_ (.A1(_02530_),
    .A2(_02538_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09653_ (.A1(_02514_),
    .A2(_02539_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09654_ (.A1(_02459_),
    .A2(_02463_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09655_ (.A1(_02456_),
    .A2(_02464_),
    .B(_02541_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09656_ (.A1(_02441_),
    .A2(_02444_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09657_ (.A1(_02441_),
    .A2(_02444_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09658_ (.A1(_02438_),
    .A2(_02543_),
    .B(_02544_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09659_ (.A1(_00373_),
    .A2(_06701_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09660_ (.A1(_00379_),
    .A2(_06691_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09661_ (.A1(_00376_),
    .A2(_06696_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09662_ (.A1(_02547_),
    .A2(_02548_),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09663_ (.A1(_02546_),
    .A2(_02549_),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09664_ (.A1(_02461_),
    .A2(_02462_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09665_ (.A1(_02461_),
    .A2(_02462_),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09666_ (.A1(_02460_),
    .A2(_02551_),
    .B(_02552_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09667_ (.A1(_00382_),
    .A2(_06685_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09668_ (.A1(_00388_),
    .A2(_06674_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09669_ (.A1(_00385_),
    .A2(_06679_),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09670_ (.A1(_02554_),
    .A2(_02555_),
    .A3(_02556_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09671_ (.A1(_02553_),
    .A2(_02557_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09672_ (.A1(_02550_),
    .A2(_02558_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09673_ (.A1(_02542_),
    .A2(_02545_),
    .A3(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09674_ (.A1(_02540_),
    .A2(_02560_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09675_ (.A1(_02512_),
    .A2(_02561_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09676_ (.A1(_02451_),
    .A2(_02465_),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09677_ (.A1(_02448_),
    .A2(_02466_),
    .B(_02563_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09678_ (.A1(_00373_),
    .A2(_06696_),
    .A3(_02455_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09679_ (.A1(_02453_),
    .A2(_02454_),
    .B(_02565_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09680_ (.A1(_02564_),
    .A2(_02566_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09681_ (.A1(_00370_),
    .A2(_06708_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09682_ (.A1(_02567_),
    .A2(_02568_),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09683_ (.A1(_02562_),
    .A2(_02569_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09684_ (.A1(_02506_),
    .A2(_02509_),
    .A3(_02570_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09685_ (.A1(_02502_),
    .A2(_02503_),
    .B(_02571_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09686_ (.A1(_02502_),
    .A2(_02503_),
    .A3(_02571_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09687_ (.A1(_02572_),
    .A2(_02573_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09688_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-11] ),
    .A2(_02501_),
    .A3(_02574_),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09689_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-12] ),
    .A2(_02495_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09690_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-13] ),
    .A2(_02394_),
    .B1(_02495_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-12] ),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09691_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-13] ),
    .A2(_02319_),
    .A3(_02393_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09692_ (.A1(_02578_),
    .A2(_02496_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09693_ (.A1(_02576_),
    .A2(_02577_),
    .B1(_02579_),
    .B2(_02405_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09694_ (.A1(_02575_),
    .A2(_02580_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09695_ (.A1(_02575_),
    .A2(_02580_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09696_ (.A1(_05182_),
    .A2(_02582_),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _09697_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[15] ),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09698_ (.A1(_05280_),
    .A2(net135),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09699_ (.A1(_02581_),
    .A2(_02583_),
    .B(_02585_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _09700_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[16] ),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09701_ (.I(_02564_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09702_ (.A1(_02587_),
    .A2(_02566_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09703_ (.A1(_02567_),
    .A2(_02568_),
    .B(_02588_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09704_ (.A1(_02512_),
    .A2(_02561_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09705_ (.A1(_02562_),
    .A2(_02569_),
    .B(_02590_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09706_ (.A1(_02513_),
    .A2(_02510_),
    .B(_02539_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09707_ (.A1(_02540_),
    .A2(_02560_),
    .B(_02592_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09708_ (.A1(_02516_),
    .A2(_02529_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09709_ (.A1(_02530_),
    .A2(_02538_),
    .B(_02594_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09710_ (.A1(_02519_),
    .A2(_02523_),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09711_ (.A1(_02524_),
    .A2(_02528_),
    .B(_02596_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09712_ (.A1(net91),
    .A2(_06710_),
    .B1(_06724_),
    .B2(net143),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09713_ (.A1(net91),
    .A2(net143),
    .A3(_06710_),
    .A4(_06724_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09714_ (.A1(_02520_),
    .A2(_02598_),
    .B(_02599_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09715_ (.A1(_00357_),
    .A2(_06738_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09716_ (.A1(_00367_),
    .A2(_06724_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09717_ (.A1(_00363_),
    .A2(_06730_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09718_ (.A1(_02601_),
    .A2(_02602_),
    .A3(_02603_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09719_ (.A1(_02600_),
    .A2(_02604_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09720_ (.A1(net96),
    .A2(_06674_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _09721_ (.A1(_00352_),
    .A2(_06744_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _09722_ (.I(_02607_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09723_ (.A1(_00355_),
    .A2(_06742_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09724_ (.A1(_02606_),
    .A2(_02608_),
    .A3(_02609_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09725_ (.A1(_02610_),
    .A2(_02605_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09726_ (.A1(_02597_),
    .A2(_02611_),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09727_ (.A1(_02526_),
    .A2(_02527_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09728_ (.A1(_02526_),
    .A2(_02527_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09729_ (.A1(_02525_),
    .A2(_02613_),
    .B(_02614_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09730_ (.A1(_06664_),
    .A2(_00398_),
    .B1(_00394_),
    .B2(_06672_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09731_ (.A1(_06664_),
    .A2(_00398_),
    .A3(_00394_),
    .A4(_06672_),
    .Z(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09732_ (.A1(_02616_),
    .A2(_02617_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09733_ (.A1(_02615_),
    .A2(_02618_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09734_ (.A1(_02535_),
    .A2(_02619_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09735_ (.A1(_02595_),
    .A2(_02612_),
    .A3(_02620_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09736_ (.I(_02557_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09737_ (.A1(_02553_),
    .A2(_02622_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09738_ (.A1(_02550_),
    .A2(_02558_),
    .B(_02623_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09739_ (.A1(_02533_),
    .A2(_02536_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09740_ (.A1(_02443_),
    .A2(_02537_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09741_ (.A1(_02625_),
    .A2(_02626_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09742_ (.A1(_00373_),
    .A2(_06708_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09743_ (.A1(_00379_),
    .A2(_06696_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09744_ (.A1(_00376_),
    .A2(_06701_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09745_ (.A1(_02629_),
    .A2(_02630_),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09746_ (.A1(_02628_),
    .A2(_02631_),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09747_ (.A1(_02555_),
    .A2(_02556_),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09748_ (.A1(_02555_),
    .A2(_02556_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09749_ (.A1(_02554_),
    .A2(_02633_),
    .B(_02634_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09750_ (.A1(_00382_),
    .A2(_06691_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09751_ (.A1(_00388_),
    .A2(_06679_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09752_ (.A1(_00385_),
    .A2(_06685_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09753_ (.A1(_02636_),
    .A2(_02637_),
    .A3(_02638_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09754_ (.A1(_02635_),
    .A2(_02639_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09755_ (.A1(_02632_),
    .A2(_02640_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09756_ (.A1(_02624_),
    .A2(_02627_),
    .A3(_02641_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09757_ (.A1(_02621_),
    .A2(_02642_),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09758_ (.A1(_02593_),
    .A2(_02643_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09759_ (.A1(_02545_),
    .A2(_02559_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09760_ (.A1(_02545_),
    .A2(_02559_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09761_ (.A1(_02542_),
    .A2(_02645_),
    .B(_02646_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09762_ (.A1(_00373_),
    .A2(_06701_),
    .A3(_02549_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09763_ (.A1(_02547_),
    .A2(_02548_),
    .B(_02648_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09764_ (.A1(_02647_),
    .A2(_02649_),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09765_ (.A1(_00370_),
    .A2(_06710_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09766_ (.A1(_02650_),
    .A2(_02651_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09767_ (.A1(_02591_),
    .A2(_02644_),
    .A3(_02652_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09768_ (.A1(_02589_),
    .A2(_02653_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09769_ (.A1(_02509_),
    .A2(_02570_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09770_ (.A1(_02509_),
    .A2(_02570_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09771_ (.A1(_02506_),
    .A2(_02655_),
    .A3(_02656_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09772_ (.A1(_02655_),
    .A2(_02657_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09773_ (.A1(_02654_),
    .A2(_02658_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09774_ (.A1(_02479_),
    .A2(_02483_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09775_ (.A1(_02660_),
    .A2(_02574_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09776_ (.I(_02572_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09777_ (.A1(_02484_),
    .A2(_02662_),
    .B(_02573_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09778_ (.I(_02663_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09779_ (.A1(_02494_),
    .A2(_02661_),
    .B(_02664_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09780_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-10] ),
    .A2(_02659_),
    .A3(_02665_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09781_ (.A1(_02501_),
    .A2(_02574_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09782_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-11] ),
    .A2(_02667_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09783_ (.A1(_02668_),
    .A2(_02582_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09784_ (.A1(_02666_),
    .A2(_02669_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09785_ (.I0(_02586_),
    .I1(_02670_),
    .S(_00395_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09786_ (.I(_02671_),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09787_ (.A1(_02578_),
    .A2(_02496_),
    .A3(_02575_),
    .A4(_02666_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09788_ (.A1(_02399_),
    .A2(_02403_),
    .B(_02672_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09789_ (.A1(_02048_),
    .A2(_02145_),
    .A3(_02397_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09790_ (.A1(_01959_),
    .A2(_01966_),
    .B(_02674_),
    .C(_02672_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09791_ (.A1(_02575_),
    .A2(_02666_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09792_ (.A1(_02659_),
    .A2(_02665_),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09793_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-11] ),
    .A2(_02667_),
    .B1(_02677_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-10] ),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09794_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-10] ),
    .A2(_02677_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _09795_ (.A1(_02576_),
    .A2(_02577_),
    .A3(_02676_),
    .B1(_02678_),
    .B2(_02679_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _09796_ (.A1(_02673_),
    .A2(_02675_),
    .A3(_02680_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09797_ (.I(_02647_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09798_ (.A1(_02682_),
    .A2(_02649_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09799_ (.A1(_02650_),
    .A2(_02651_),
    .B(_02683_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09800_ (.A1(_02593_),
    .A2(_02643_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09801_ (.A1(_02644_),
    .A2(_02652_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09802_ (.A1(_02685_),
    .A2(_02686_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09803_ (.A1(_02620_),
    .A2(_02612_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09804_ (.A1(_02612_),
    .A2(_02620_),
    .ZN(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09805_ (.A1(_02595_),
    .A2(_02688_),
    .A3(_02689_),
    .B1(_02621_),
    .B2(_02642_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09806_ (.A1(net151),
    .A2(_02611_),
    .B(_02688_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09807_ (.A1(net150),
    .A2(_02604_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09808_ (.A1(_02605_),
    .A2(net149),
    .B(_02692_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09809_ (.A1(net61),
    .A2(_06724_),
    .B1(_06730_),
    .B2(net60),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09810_ (.A1(net61),
    .A2(net60),
    .A3(_06724_),
    .A4(_06730_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09811_ (.A1(_02601_),
    .A2(_02694_),
    .B(_02695_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09812_ (.A1(net73),
    .A2(_06742_),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09813_ (.A1(net91),
    .A2(_06730_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09814_ (.A1(net60),
    .A2(_06738_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09815_ (.A1(_02697_),
    .A2(_02698_),
    .A3(_02699_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09816_ (.A1(_02696_),
    .A2(_02700_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09817_ (.A1(net95),
    .A2(_06679_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09818_ (.A1(_00355_),
    .A2(_06744_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _09819_ (.I(_02703_),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09820_ (.A1(_02608_),
    .A2(_02702_),
    .A3(_02704_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09821_ (.A1(_02701_),
    .A2(_02705_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09822_ (.A1(_02693_),
    .A2(_02706_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09823_ (.A1(net63),
    .A2(_06674_),
    .B(_02608_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09824_ (.A1(net63),
    .A2(_06674_),
    .A3(_02608_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09825_ (.A1(_02708_),
    .A2(_02609_),
    .B(_02709_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09826_ (.A1(_00398_),
    .A2(_06672_),
    .B1(_06674_),
    .B2(_00394_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09827_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06672_),
    .A4(_06674_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09828_ (.A1(_02711_),
    .A2(_02712_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09829_ (.A1(_02710_),
    .A2(_02713_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09830_ (.A1(_02617_),
    .A2(_02714_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09831_ (.A1(_02691_),
    .A2(_02707_),
    .A3(_02715_),
    .Z(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09832_ (.A1(_02635_),
    .A2(_02639_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09833_ (.A1(_02632_),
    .A2(_02640_),
    .B(_02717_),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09834_ (.A1(_02615_),
    .A2(_02618_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09835_ (.A1(_02535_),
    .A2(_02619_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09836_ (.A1(_02719_),
    .A2(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09837_ (.A1(_00373_),
    .A2(_06710_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09838_ (.A1(_00379_),
    .A2(_06701_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09839_ (.A1(_00376_),
    .A2(_06708_),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09840_ (.A1(_02723_),
    .A2(_02724_),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09841_ (.A1(_02722_),
    .A2(_02725_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09842_ (.A1(_02637_),
    .A2(_02638_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09843_ (.A1(_02637_),
    .A2(_02638_),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09844_ (.A1(_02636_),
    .A2(_02727_),
    .B(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09845_ (.A1(_00382_),
    .A2(_06696_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09846_ (.A1(_00388_),
    .A2(_06685_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09847_ (.A1(_00385_),
    .A2(_06691_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09848_ (.A1(_02730_),
    .A2(_02731_),
    .A3(_02732_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09849_ (.A1(_02729_),
    .A2(_02733_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09850_ (.A1(_02726_),
    .A2(_02734_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09851_ (.A1(_02718_),
    .A2(_02721_),
    .A3(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09852_ (.A1(_02736_),
    .A2(_02716_),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09853_ (.A1(_02690_),
    .A2(_02737_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09854_ (.A1(_02627_),
    .A2(_02641_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09855_ (.A1(_02627_),
    .A2(_02641_),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09856_ (.A1(_02624_),
    .A2(_02739_),
    .B(_02740_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09857_ (.A1(_00373_),
    .A2(_06708_),
    .A3(_02631_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09858_ (.A1(_02629_),
    .A2(_02630_),
    .B(_02742_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09859_ (.A1(_02741_),
    .A2(_02743_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09860_ (.A1(_00370_),
    .A2(_06724_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09861_ (.A1(_02744_),
    .A2(_02745_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09862_ (.A1(_02746_),
    .A2(_02738_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09863_ (.A1(_02687_),
    .A2(_02747_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09864_ (.A1(_02684_),
    .A2(_02748_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09865_ (.A1(_02644_),
    .A2(_02652_),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09866_ (.A1(_02644_),
    .A2(_02652_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09867_ (.A1(_02589_),
    .A2(_02653_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09868_ (.A1(_02591_),
    .A2(_02750_),
    .A3(_02751_),
    .B(_02752_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09869_ (.A1(_02749_),
    .A2(_02753_),
    .Z(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09870_ (.I(_02754_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09871_ (.A1(_02654_),
    .A2(_02658_),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09872_ (.A1(_02659_),
    .A2(_02665_),
    .B(_02756_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09873_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ),
    .A2(_02755_),
    .A3(_02757_),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09874_ (.I(_02758_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09875_ (.A1(_02681_),
    .A2(_02759_),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09876_ (.A1(_02681_),
    .A2(_02759_),
    .B(_05182_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _09877_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[17] ),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09878_ (.A1(_05280_),
    .A2(_02762_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09879_ (.A1(_02760_),
    .A2(_02761_),
    .B(_02763_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09880_ (.I(_02741_),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09881_ (.A1(_02764_),
    .A2(_02743_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09882_ (.A1(_02744_),
    .A2(_02745_),
    .B(_02765_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09883_ (.A1(_02690_),
    .A2(_02737_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09884_ (.A1(_02738_),
    .A2(_02746_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09885_ (.A1(_02767_),
    .A2(_02768_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09886_ (.A1(_02707_),
    .A2(_02715_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09887_ (.A1(_02707_),
    .A2(_02715_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09888_ (.A1(_02691_),
    .A2(_02770_),
    .A3(_02771_),
    .B1(_02716_),
    .B2(_02736_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09889_ (.A1(_02693_),
    .A2(_02706_),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09890_ (.A1(_02696_),
    .A2(_02700_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09891_ (.A1(_02701_),
    .A2(_02705_),
    .B(_02774_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09892_ (.A1(net61),
    .A2(_06730_),
    .B1(_06738_),
    .B2(net60),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09893_ (.A1(net61),
    .A2(net60),
    .A3(_06730_),
    .A4(_06738_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09894_ (.A1(_02697_),
    .A2(_02776_),
    .B(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09895_ (.A1(net73),
    .A2(_06744_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09896_ (.A1(net61),
    .A2(_06738_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09897_ (.A1(net60),
    .A2(_06742_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09898_ (.A1(_02779_),
    .A2(_02780_),
    .A3(_02781_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09899_ (.A1(_02778_),
    .A2(_02782_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09900_ (.A1(net95),
    .A2(_06685_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09901_ (.A1(_02608_),
    .A2(_02704_),
    .A3(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09902_ (.A1(_02783_),
    .A2(_02785_),
    .Z(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09903_ (.A1(_02775_),
    .A2(_02786_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09904_ (.A1(net63),
    .A2(_06679_),
    .B(_02608_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09905_ (.A1(net63),
    .A2(_06679_),
    .A3(_02608_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09906_ (.A1(_02788_),
    .A2(_02704_),
    .B(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09907_ (.A1(_00398_),
    .A2(_06674_),
    .B1(_06679_),
    .B2(_00394_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09908_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06674_),
    .A4(_06679_),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09909_ (.A1(_02791_),
    .A2(_02792_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09910_ (.A1(_02790_),
    .A2(_02793_),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09911_ (.A1(_02712_),
    .A2(_02794_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09912_ (.A1(_02787_),
    .A2(_02795_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09913_ (.A1(_02773_),
    .A2(_02770_),
    .B(_02796_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09914_ (.A1(_02773_),
    .A2(_02770_),
    .A3(_02796_),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09915_ (.A1(_02797_),
    .A2(_02798_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09916_ (.A1(_02729_),
    .A2(_02733_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09917_ (.A1(_02726_),
    .A2(_02734_),
    .B(_02800_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09918_ (.A1(_02710_),
    .A2(_02713_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09919_ (.A1(_02617_),
    .A2(_02714_),
    .B(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09920_ (.A1(_00373_),
    .A2(_06724_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09921_ (.A1(_00379_),
    .A2(_06708_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09922_ (.A1(_00376_),
    .A2(_06710_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09923_ (.A1(_02805_),
    .A2(_02806_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09924_ (.A1(_02804_),
    .A2(_02807_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09925_ (.A1(_02731_),
    .A2(_02732_),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09926_ (.A1(_02731_),
    .A2(_02732_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09927_ (.A1(_02730_),
    .A2(_02809_),
    .B(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09928_ (.A1(_00382_),
    .A2(_06701_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09929_ (.A1(_00388_),
    .A2(_00385_),
    .A3(_06691_),
    .A4(_06696_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09930_ (.A1(_00388_),
    .A2(_06691_),
    .B1(_06696_),
    .B2(_00385_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09931_ (.A1(_02812_),
    .A2(_02813_),
    .A3(_02814_),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09932_ (.A1(_02813_),
    .A2(_02814_),
    .B(_02812_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09933_ (.A1(_02815_),
    .A2(_02816_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09934_ (.A1(_02811_),
    .A2(_02817_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09935_ (.A1(_02808_),
    .A2(_02818_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09936_ (.A1(_02801_),
    .A2(_02803_),
    .A3(_02819_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09937_ (.A1(_02799_),
    .A2(_02820_),
    .Z(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09938_ (.A1(_02772_),
    .A2(_02821_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09939_ (.A1(_02721_),
    .A2(_02735_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09940_ (.A1(_02721_),
    .A2(_02735_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09941_ (.A1(_02718_),
    .A2(_02823_),
    .B(_02824_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09942_ (.I(_02825_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09943_ (.A1(_00373_),
    .A2(_06710_),
    .A3(_02725_),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09944_ (.A1(_02723_),
    .A2(_02724_),
    .B(_02827_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09945_ (.A1(_02826_),
    .A2(_02828_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09946_ (.A1(_00370_),
    .A2(_06730_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09947_ (.A1(_02829_),
    .A2(_02830_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09948_ (.A1(_02822_),
    .A2(_02831_),
    .Z(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09949_ (.A1(_02769_),
    .A2(_02832_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09950_ (.A1(_02766_),
    .A2(_02833_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09951_ (.A1(_02687_),
    .A2(_02747_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09952_ (.A1(_02684_),
    .A2(_02748_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09953_ (.A1(_02835_),
    .A2(_02836_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09954_ (.A1(_02834_),
    .A2(_02837_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09955_ (.A1(_02660_),
    .A2(_02574_),
    .A3(_02659_),
    .A4(_02755_),
    .Z(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09956_ (.A1(_02493_),
    .A2(_02839_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09957_ (.I(_02749_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09958_ (.A1(_02841_),
    .A2(_02753_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09959_ (.A1(_02659_),
    .A2(_02663_),
    .A3(_02755_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09960_ (.A1(_02841_),
    .A2(_02753_),
    .B(_02756_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09961_ (.A1(_02842_),
    .A2(_02843_),
    .A3(_02844_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09962_ (.A1(net55),
    .A2(_02839_),
    .B(_02840_),
    .C(_02845_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09963_ (.A1(_02838_),
    .A2(_02846_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09964_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-8] ),
    .A2(_02847_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09965_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-8] ),
    .A2(_02847_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09966_ (.A1(_02848_),
    .A2(_02849_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09967_ (.A1(net53),
    .A2(_02757_),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09968_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ),
    .A2(_02851_),
    .B(_02760_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09969_ (.A1(_02850_),
    .A2(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _09970_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[18] ),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09971_ (.A1(_05280_),
    .A2(_02854_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09972_ (.A1(_05822_),
    .A2(_02853_),
    .B(_02855_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09973_ (.A1(_02769_),
    .A2(_02832_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09974_ (.A1(_02766_),
    .A2(_02833_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09975_ (.A1(_02826_),
    .A2(_02828_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09976_ (.A1(_00370_),
    .A2(_06730_),
    .A3(_02829_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09977_ (.A1(_02858_),
    .A2(_02859_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09978_ (.A1(_02772_),
    .A2(_02821_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09979_ (.A1(_02822_),
    .A2(_02831_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09980_ (.A1(_02861_),
    .A2(_02862_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09981_ (.A1(_02799_),
    .A2(_02820_),
    .B(_02797_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09982_ (.A1(_02775_),
    .A2(_02786_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09983_ (.A1(_02787_),
    .A2(_02795_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09984_ (.A1(_02865_),
    .A2(_02866_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09985_ (.A1(_02778_),
    .A2(_02782_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09986_ (.A1(_02783_),
    .A2(_02785_),
    .B(_02868_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09987_ (.A1(net61),
    .A2(_06738_),
    .B1(_06742_),
    .B2(net60),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09988_ (.A1(net61),
    .A2(net60),
    .A3(_06738_),
    .A4(_06742_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09989_ (.A1(_02779_),
    .A2(_02870_),
    .B(_02871_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09990_ (.A1(net61),
    .A2(_06742_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09991_ (.A1(net60),
    .A2(_06744_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09992_ (.A1(_02779_),
    .A2(_02873_),
    .A3(_02874_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09993_ (.A1(_02872_),
    .A2(_02875_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09994_ (.A1(net63),
    .A2(_06691_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09995_ (.A1(_02608_),
    .A2(_02704_),
    .A3(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09996_ (.A1(_02876_),
    .A2(_02878_),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09997_ (.A1(_02869_),
    .A2(_02879_),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09998_ (.A1(net63),
    .A2(_06685_),
    .B(_02608_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09999_ (.A1(net63),
    .A2(_06685_),
    .A3(_02608_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10000_ (.A1(_02704_),
    .A2(_02881_),
    .B(_02882_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10001_ (.A1(_00398_),
    .A2(_06679_),
    .B1(_06685_),
    .B2(_00394_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10002_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06679_),
    .A4(_06685_),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10003_ (.A1(_02884_),
    .A2(_02885_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10004_ (.A1(_02883_),
    .A2(_02886_),
    .Z(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10005_ (.A1(_02792_),
    .A2(_02887_),
    .Z(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10006_ (.A1(_02880_),
    .A2(_02888_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10007_ (.A1(_02867_),
    .A2(_02889_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10008_ (.A1(_02811_),
    .A2(_02815_),
    .A3(_02816_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10009_ (.A1(_02808_),
    .A2(_02818_),
    .B(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10010_ (.A1(_02790_),
    .A2(_02793_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10011_ (.A1(_02712_),
    .A2(_02794_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10012_ (.A1(_02893_),
    .A2(_02894_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10013_ (.A1(_00373_),
    .A2(_06730_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10014_ (.A1(_00379_),
    .A2(_06710_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10015_ (.A1(_00376_),
    .A2(_06724_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10016_ (.A1(_02897_),
    .A2(_02898_),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10017_ (.A1(_02896_),
    .A2(_02899_),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10018_ (.A1(_02812_),
    .A2(_02813_),
    .A3(_02814_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10019_ (.A1(_02813_),
    .A2(_02901_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10020_ (.A1(_00382_),
    .A2(_06708_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10021_ (.A1(_00388_),
    .A2(_06696_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10022_ (.A1(_00385_),
    .A2(_06701_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10023_ (.A1(_02903_),
    .A2(_02904_),
    .A3(_02905_),
    .Z(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10024_ (.A1(_02902_),
    .A2(_02906_),
    .Z(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10025_ (.A1(_02902_),
    .A2(_02906_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10026_ (.A1(_02907_),
    .A2(_02908_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10027_ (.A1(_02900_),
    .A2(_02909_),
    .Z(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10028_ (.A1(_02892_),
    .A2(_02895_),
    .A3(_02910_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10029_ (.A1(_02890_),
    .A2(_02911_),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10030_ (.A1(_02864_),
    .A2(_02912_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10031_ (.A1(_02803_),
    .A2(_02819_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10032_ (.A1(_02803_),
    .A2(_02819_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10033_ (.A1(_02801_),
    .A2(_02914_),
    .B(_02915_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10034_ (.A1(_00373_),
    .A2(_06724_),
    .A3(_02807_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10035_ (.A1(_02805_),
    .A2(_02806_),
    .B(_02917_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10036_ (.A1(_02916_),
    .A2(_02918_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10037_ (.A1(_00370_),
    .A2(_06738_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10038_ (.A1(_02919_),
    .A2(_02920_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10039_ (.A1(_02913_),
    .A2(_02921_),
    .Z(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10040_ (.A1(_02860_),
    .A2(_02863_),
    .A3(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10041_ (.A1(_02856_),
    .A2(_02857_),
    .B(_02923_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10042_ (.A1(_02856_),
    .A2(_02857_),
    .A3(_02923_),
    .Z(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10043_ (.A1(_02924_),
    .A2(_02925_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10044_ (.A1(_02834_),
    .A2(_02837_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10045_ (.A1(_02838_),
    .A2(_02846_),
    .B(_02927_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10046_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-7] ),
    .A2(_02926_),
    .A3(_02928_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10047_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ),
    .A2(_02851_),
    .B(_02848_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10048_ (.A1(_02849_),
    .A2(_02930_),
    .Z(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10049_ (.A1(_02758_),
    .A2(_02850_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10050_ (.A1(_02681_),
    .A2(_02932_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10051_ (.A1(_02931_),
    .A2(_02933_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10052_ (.A1(_02929_),
    .A2(_02934_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10053_ (.A1(_02929_),
    .A2(_02934_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10054_ (.A1(_05182_),
    .A2(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10055_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[19] ),
    .Z(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10056_ (.A1(_05280_),
    .A2(_02938_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10057_ (.A1(_02935_),
    .A2(_02937_),
    .B(_02939_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10058_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[20] ),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10059_ (.I(_02916_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10060_ (.A1(_02941_),
    .A2(_02918_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10061_ (.A1(_02919_),
    .A2(_02920_),
    .B(_02942_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10062_ (.A1(_02864_),
    .A2(_02912_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10063_ (.A1(_02913_),
    .A2(_02921_),
    .B(_02944_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10064_ (.A1(_02867_),
    .A2(_02889_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10065_ (.A1(_02890_),
    .A2(_02911_),
    .B(_02946_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10066_ (.A1(_02869_),
    .A2(_02879_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10067_ (.A1(_02880_),
    .A2(_02888_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10068_ (.A1(_02948_),
    .A2(_02949_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10069_ (.A1(_02872_),
    .A2(_02875_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10070_ (.A1(_02876_),
    .A2(_02878_),
    .B(_02951_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10071_ (.A1(net95),
    .A2(_06696_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10072_ (.A1(_02608_),
    .A2(_02704_),
    .A3(_02953_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10073_ (.A1(net61),
    .A2(_06744_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10074_ (.A1(_02873_),
    .A2(_02874_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10075_ (.A1(_02873_),
    .A2(_02874_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10076_ (.A1(net161),
    .A2(_02956_),
    .B1(_02957_),
    .B2(_02779_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10077_ (.A1(_02874_),
    .A2(_02955_),
    .A3(_02958_),
    .Z(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10078_ (.A1(_02954_),
    .A2(_02959_),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10079_ (.A1(_02952_),
    .A2(_02960_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10080_ (.A1(net63),
    .A2(_06691_),
    .B(_02608_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10081_ (.A1(net63),
    .A2(_06691_),
    .A3(_02608_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10082_ (.A1(_02704_),
    .A2(_02962_),
    .B(_02963_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10083_ (.A1(_00398_),
    .A2(_06685_),
    .B1(_06691_),
    .B2(_00394_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10084_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06685_),
    .A4(_06691_),
    .Z(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10085_ (.A1(_02965_),
    .A2(_02966_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10086_ (.A1(_02964_),
    .A2(_02967_),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10087_ (.A1(_02885_),
    .A2(_02968_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10088_ (.A1(_02961_),
    .A2(_02969_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10089_ (.A1(_02950_),
    .A2(_02970_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10090_ (.A1(_02900_),
    .A2(_02909_),
    .B(_02907_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10091_ (.A1(_02883_),
    .A2(_02886_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10092_ (.A1(_02792_),
    .A2(_02887_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10093_ (.A1(_02973_),
    .A2(_02974_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10094_ (.A1(_00373_),
    .A2(_06738_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10095_ (.A1(_00379_),
    .A2(_06724_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10096_ (.A1(_00376_),
    .A2(_06730_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10097_ (.A1(_02977_),
    .A2(_02978_),
    .Z(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10098_ (.A1(_02976_),
    .A2(_02979_),
    .Z(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10099_ (.A1(_02904_),
    .A2(_02905_),
    .Z(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10100_ (.A1(_02904_),
    .A2(_02905_),
    .Z(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10101_ (.A1(_02903_),
    .A2(_02981_),
    .B(_02982_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10102_ (.A1(_00382_),
    .A2(_06710_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10103_ (.A1(_00388_),
    .A2(_06701_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10104_ (.A1(_00385_),
    .A2(_06708_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10105_ (.A1(_02984_),
    .A2(_02985_),
    .A3(_02986_),
    .Z(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10106_ (.A1(_02983_),
    .A2(_02987_),
    .Z(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10107_ (.A1(_02980_),
    .A2(_02988_),
    .Z(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10108_ (.A1(_02972_),
    .A2(_02975_),
    .A3(_02989_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10109_ (.A1(_02971_),
    .A2(_02990_),
    .Z(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10110_ (.A1(_02947_),
    .A2(_02991_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10111_ (.A1(_02895_),
    .A2(_02910_),
    .Z(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10112_ (.A1(_02895_),
    .A2(_02910_),
    .Z(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10113_ (.A1(_02892_),
    .A2(_02993_),
    .B(_02994_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10114_ (.A1(_00373_),
    .A2(_06730_),
    .A3(_02899_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10115_ (.A1(_02897_),
    .A2(_02898_),
    .B(_02996_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10116_ (.A1(_02995_),
    .A2(_02997_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10117_ (.A1(_00370_),
    .A2(_06742_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10118_ (.A1(_02998_),
    .A2(_02999_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10119_ (.A1(_02992_),
    .A2(_03000_),
    .Z(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10120_ (.A1(_02945_),
    .A2(_03001_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10121_ (.A1(_02943_),
    .A2(_03002_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10122_ (.A1(_02863_),
    .A2(_02922_),
    .Z(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10123_ (.A1(_02863_),
    .A2(_02922_),
    .Z(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10124_ (.A1(_02860_),
    .A2(_03004_),
    .B(_03005_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10125_ (.A1(_03003_),
    .A2(_03006_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10126_ (.I(_02838_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10127_ (.A1(_03008_),
    .A2(_02926_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10128_ (.A1(_02834_),
    .A2(_02837_),
    .B(_02924_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10129_ (.A1(_02925_),
    .A2(_03010_),
    .Z(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10130_ (.A1(_02846_),
    .A2(_03009_),
    .B(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10131_ (.A1(_00506_),
    .A2(_03007_),
    .A3(_03012_),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10132_ (.A1(_02926_),
    .A2(_02928_),
    .Z(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10133_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-7] ),
    .A2(_03014_),
    .B(_02935_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10134_ (.A1(_03013_),
    .A2(_03015_),
    .Z(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10135_ (.I0(_02940_),
    .I1(_03016_),
    .S(_00395_),
    .Z(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10136_ (.I(_03017_),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10137_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[21] ),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10138_ (.A1(_05822_),
    .A2(_03018_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10139_ (.I(_02995_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10140_ (.A1(_03020_),
    .A2(_02997_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10141_ (.A1(_02998_),
    .A2(_02999_),
    .B(_03021_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10142_ (.A1(_02947_),
    .A2(_02991_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10143_ (.A1(_02992_),
    .A2(_03000_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10144_ (.A1(_03023_),
    .A2(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10145_ (.A1(_02950_),
    .A2(_02970_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10146_ (.A1(_02971_),
    .A2(_02990_),
    .B(_03026_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10147_ (.A1(_02952_),
    .A2(_02960_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10148_ (.A1(_02961_),
    .A2(_02969_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10149_ (.A1(_03028_),
    .A2(_03029_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10150_ (.A1(_00358_),
    .A2(_02874_),
    .A3(_02955_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10151_ (.A1(_02954_),
    .A2(_02959_),
    .B(_03031_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10152_ (.A1(net63),
    .A2(_06701_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10153_ (.A1(_02608_),
    .A2(_02704_),
    .A3(_03033_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10154_ (.A1(net61),
    .A2(net60),
    .B(_06744_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10155_ (.A1(_02779_),
    .A2(_03035_),
    .B(_03031_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10156_ (.I(_03036_),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10157_ (.A1(_03034_),
    .A2(_03037_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10158_ (.A1(_03032_),
    .A2(_03038_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10159_ (.A1(net63),
    .A2(_06696_),
    .B(_02608_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10160_ (.A1(net63),
    .A2(_06696_),
    .A3(_02608_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10161_ (.A1(_02704_),
    .A2(_03040_),
    .B(_03041_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10162_ (.A1(_00398_),
    .A2(_06691_),
    .B1(_06696_),
    .B2(_00394_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10163_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06691_),
    .A4(_06696_),
    .Z(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10164_ (.A1(_03043_),
    .A2(_03044_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10165_ (.A1(_03042_),
    .A2(_03045_),
    .Z(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10166_ (.A1(_02966_),
    .A2(_03046_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10167_ (.A1(_03039_),
    .A2(_03047_),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10168_ (.A1(_03030_),
    .A2(_03048_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10169_ (.I(_02987_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10170_ (.A1(_02983_),
    .A2(_03050_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10171_ (.A1(_02980_),
    .A2(_02988_),
    .B(_03051_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10172_ (.A1(_02964_),
    .A2(_02967_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10173_ (.A1(_02885_),
    .A2(_02968_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10174_ (.A1(_03053_),
    .A2(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10175_ (.A1(_00373_),
    .A2(_06742_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10176_ (.A1(_00379_),
    .A2(_06730_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10177_ (.A1(_00376_),
    .A2(_06738_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10178_ (.A1(_03057_),
    .A2(_03058_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10179_ (.A1(_03056_),
    .A2(_03059_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10180_ (.A1(_02985_),
    .A2(_02986_),
    .Z(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10181_ (.A1(_02985_),
    .A2(_02986_),
    .Z(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10182_ (.A1(_02984_),
    .A2(_03061_),
    .B(_03062_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10183_ (.A1(_00382_),
    .A2(_06724_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10184_ (.A1(_00388_),
    .A2(_06708_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10185_ (.A1(_00385_),
    .A2(_06710_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10186_ (.A1(_03064_),
    .A2(_03065_),
    .A3(_03066_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10187_ (.A1(_03063_),
    .A2(_03067_),
    .Z(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10188_ (.A1(_03060_),
    .A2(_03068_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10189_ (.A1(_03052_),
    .A2(_03055_),
    .A3(_03069_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10190_ (.A1(_03049_),
    .A2(_03070_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10191_ (.A1(_03027_),
    .A2(_03071_),
    .Z(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10192_ (.A1(_02977_),
    .A2(_02978_),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10193_ (.A1(_00373_),
    .A2(_06738_),
    .A3(_02979_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10194_ (.A1(_02975_),
    .A2(_02989_),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10195_ (.A1(_02975_),
    .A2(_02989_),
    .Z(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10196_ (.A1(_02972_),
    .A2(_03075_),
    .B(_03076_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10197_ (.A1(_03073_),
    .A2(_03074_),
    .B(_03077_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10198_ (.A1(_03073_),
    .A2(_03074_),
    .A3(_03077_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10199_ (.A1(_03078_),
    .A2(_03079_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10200_ (.A1(_00370_),
    .A2(_06744_),
    .Z(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10201_ (.I(_03081_),
    .Z(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10202_ (.A1(_03080_),
    .A2(_03082_),
    .Z(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10203_ (.A1(_03072_),
    .A2(_03083_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10204_ (.A1(_03022_),
    .A2(_03025_),
    .A3(_03084_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10205_ (.I(_02945_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10206_ (.A1(_03086_),
    .A2(_03001_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10207_ (.A1(_02943_),
    .A2(_03002_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10208_ (.A1(_03087_),
    .A2(_03088_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10209_ (.A1(_03085_),
    .A2(_03089_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10210_ (.I(_03090_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10211_ (.A1(_03003_),
    .A2(_03006_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10212_ (.A1(_03007_),
    .A2(_03012_),
    .B(_03092_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10213_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ),
    .A2(_03091_),
    .A3(_03093_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10214_ (.I(_03094_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _10215_ (.A1(_02929_),
    .A2(_03013_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10216_ (.A1(_03007_),
    .A2(_03012_),
    .Z(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _10217_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-7] ),
    .A2(_03014_),
    .B1(_03097_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-6] ),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10218_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-6] ),
    .A2(_03097_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10219_ (.A1(_02758_),
    .A2(_02850_),
    .A3(_03096_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _10220_ (.A1(_02673_),
    .A2(_02675_),
    .A3(_02680_),
    .B(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _10221_ (.A1(_02931_),
    .A2(_03096_),
    .B1(_03098_),
    .B2(_03099_),
    .C(_03101_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10222_ (.A1(_03095_),
    .A2(_03102_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10223_ (.A1(_03095_),
    .A2(_03102_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10224_ (.A1(_05387_),
    .A2(_03103_),
    .A3(_03104_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10225_ (.A1(_03019_),
    .A2(_03105_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10226_ (.A1(_03080_),
    .A2(_03082_),
    .B(_03078_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10227_ (.I(_03106_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10228_ (.A1(_03027_),
    .A2(_03071_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10229_ (.A1(_03072_),
    .A2(_03083_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10230_ (.A1(_03108_),
    .A2(_03109_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10231_ (.A1(_03030_),
    .A2(_03048_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10232_ (.A1(_03049_),
    .A2(_03070_),
    .B(_03111_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10233_ (.A1(_03032_),
    .A2(_03038_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10234_ (.A1(_03039_),
    .A2(_03047_),
    .B(_03113_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10235_ (.A1(net61),
    .A2(net60),
    .A3(net161),
    .A4(_06744_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10236_ (.A1(_03034_),
    .A2(_03037_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10237_ (.A1(_03115_),
    .A2(_03116_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10238_ (.A1(net63),
    .A2(_06708_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10239_ (.A1(_02608_),
    .A2(_02704_),
    .A3(_03118_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10240_ (.A1(_03037_),
    .A2(_03119_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10241_ (.A1(_03117_),
    .A2(_03120_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10242_ (.A1(net63),
    .A2(_06701_),
    .B(net57),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10243_ (.A1(net63),
    .A2(_06701_),
    .A3(net57),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10244_ (.A1(_02704_),
    .A2(_03122_),
    .B(_03123_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10245_ (.A1(_00398_),
    .A2(_06696_),
    .B1(_06701_),
    .B2(_00394_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10246_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06696_),
    .A4(_06701_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10247_ (.A1(_03125_),
    .A2(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10248_ (.A1(_03124_),
    .A2(_03127_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10249_ (.A1(_03044_),
    .A2(_03128_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10250_ (.A1(_03121_),
    .A2(_03129_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10251_ (.A1(_03114_),
    .A2(_03130_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10252_ (.I(_03067_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10253_ (.A1(_03063_),
    .A2(_03132_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10254_ (.A1(_03060_),
    .A2(_03068_),
    .B(_03133_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10255_ (.A1(_03042_),
    .A2(_03045_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10256_ (.A1(_02966_),
    .A2(_03046_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10257_ (.A1(_03135_),
    .A2(_03136_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10258_ (.A1(_00373_),
    .A2(_06744_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10259_ (.A1(_00379_),
    .A2(_06738_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10260_ (.A1(_00376_),
    .A2(_06742_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10261_ (.A1(_03139_),
    .A2(_03140_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10262_ (.A1(_03138_),
    .A2(_03141_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10263_ (.A1(_03065_),
    .A2(_03066_),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10264_ (.A1(_03065_),
    .A2(_03066_),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10265_ (.A1(_03064_),
    .A2(_03143_),
    .B(_03144_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10266_ (.A1(_00382_),
    .A2(_06730_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10267_ (.A1(_00388_),
    .A2(_06710_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10268_ (.A1(_00385_),
    .A2(_06724_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10269_ (.A1(_03146_),
    .A2(_03147_),
    .A3(_03148_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10270_ (.A1(_03145_),
    .A2(_03149_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10271_ (.A1(_03142_),
    .A2(_03150_),
    .Z(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10272_ (.A1(_03134_),
    .A2(_03137_),
    .A3(_03151_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10273_ (.A1(_03131_),
    .A2(_03152_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10274_ (.A1(_03112_),
    .A2(_03153_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10275_ (.A1(_03057_),
    .A2(_03058_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10276_ (.A1(_00373_),
    .A2(_06742_),
    .A3(_03059_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10277_ (.A1(_03055_),
    .A2(_03069_),
    .Z(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10278_ (.A1(_03055_),
    .A2(_03069_),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10279_ (.A1(_03052_),
    .A2(_03157_),
    .B(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10280_ (.A1(_03155_),
    .A2(_03156_),
    .B(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10281_ (.A1(_03155_),
    .A2(_03156_),
    .A3(_03159_),
    .Z(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10282_ (.A1(_03160_),
    .A2(_03161_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10283_ (.A1(_03082_),
    .A2(_03162_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10284_ (.A1(_03154_),
    .A2(_03163_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10285_ (.A1(_03110_),
    .A2(_03164_),
    .Z(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10286_ (.A1(_03107_),
    .A2(_03165_),
    .Z(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10287_ (.A1(_03025_),
    .A2(_03084_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10288_ (.A1(_03025_),
    .A2(_03084_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10289_ (.A1(_03022_),
    .A2(_03167_),
    .B(_03168_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10290_ (.A1(_03166_),
    .A2(_03169_),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10291_ (.I(_03085_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10292_ (.A1(_03007_),
    .A2(_03091_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10293_ (.A1(_03009_),
    .A2(_03172_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10294_ (.A1(_02225_),
    .A2(_02226_),
    .A3(_02490_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10295_ (.A1(_02141_),
    .A2(_02142_),
    .B(_03174_),
    .C(_02140_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10296_ (.I(_02839_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10297_ (.A1(_02839_),
    .A2(_02493_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _10298_ (.A1(_02842_),
    .A2(_02843_),
    .A3(_02844_),
    .Z(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10299_ (.A1(_03175_),
    .A2(_03176_),
    .B(_03177_),
    .C(_03178_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10300_ (.A1(_03171_),
    .A2(_03089_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10301_ (.A1(_03003_),
    .A2(_03006_),
    .A3(_03180_),
    .B1(_03172_),
    .B2(_03011_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10302_ (.A1(_03171_),
    .A2(_03089_),
    .B1(_03173_),
    .B2(_03179_),
    .C(_03181_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10303_ (.A1(_03182_),
    .A2(_03170_),
    .Z(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10304_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-4] ),
    .A2(_03183_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10305_ (.A1(_03090_),
    .A2(_03093_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10306_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ),
    .A2(_03185_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10307_ (.A1(_03186_),
    .A2(_03104_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10308_ (.A1(_03184_),
    .A2(_03187_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10309_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[22] ),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10310_ (.A1(_05280_),
    .A2(_03189_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10311_ (.A1(_05822_),
    .A2(_03188_),
    .B(_03190_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10312_ (.A1(_03082_),
    .A2(_03162_),
    .B(_03160_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10313_ (.A1(_03112_),
    .A2(_03153_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10314_ (.A1(_03154_),
    .A2(_03163_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10315_ (.A1(_03192_),
    .A2(_03193_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10316_ (.A1(_03114_),
    .A2(_03130_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10317_ (.A1(_03131_),
    .A2(_03152_),
    .B(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10318_ (.A1(_03117_),
    .A2(_03120_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10319_ (.A1(_03121_),
    .A2(_03129_),
    .B(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10320_ (.A1(_03037_),
    .A2(_03119_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10321_ (.A1(_03115_),
    .A2(_03199_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10322_ (.A1(net63),
    .A2(_06710_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10323_ (.A1(_02608_),
    .A2(_02704_),
    .A3(_03201_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10324_ (.A1(_03037_),
    .A2(_03202_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10325_ (.A1(_03200_),
    .A2(_03203_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10326_ (.A1(net63),
    .A2(_06708_),
    .B(net57),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10327_ (.A1(net63),
    .A2(_06708_),
    .A3(net57),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10328_ (.A1(_02704_),
    .A2(_03205_),
    .B(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10329_ (.A1(_00398_),
    .A2(_06701_),
    .B1(_06708_),
    .B2(_00394_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10330_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06701_),
    .A4(_06708_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10331_ (.A1(_03208_),
    .A2(_03209_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10332_ (.A1(_03207_),
    .A2(_03210_),
    .Z(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10333_ (.A1(_03126_),
    .A2(_03211_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10334_ (.A1(_03204_),
    .A2(_03212_),
    .Z(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10335_ (.A1(_03198_),
    .A2(_03213_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10336_ (.I(_03149_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10337_ (.A1(_03145_),
    .A2(_03215_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10338_ (.A1(_03142_),
    .A2(_03150_),
    .B(_03216_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10339_ (.I(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10340_ (.A1(_03124_),
    .A2(_03127_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10341_ (.A1(_03044_),
    .A2(_03128_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10342_ (.A1(_03219_),
    .A2(_03220_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10343_ (.A1(_00379_),
    .A2(_06742_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10344_ (.A1(_00376_),
    .A2(_06744_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10345_ (.A1(_03222_),
    .A2(_03223_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10346_ (.A1(_03222_),
    .A2(_03223_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10347_ (.A1(_03224_),
    .A2(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10348_ (.A1(_03138_),
    .A2(_03226_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10349_ (.A1(_03147_),
    .A2(_03148_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10350_ (.A1(_03147_),
    .A2(_03148_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10351_ (.A1(_03146_),
    .A2(_03228_),
    .B(_03229_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10352_ (.A1(_00382_),
    .A2(_06738_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10353_ (.A1(_00388_),
    .A2(_06724_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10354_ (.A1(_00385_),
    .A2(_06730_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10355_ (.A1(_03231_),
    .A2(_03232_),
    .A3(_03233_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10356_ (.A1(_03230_),
    .A2(_03234_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10357_ (.A1(_03227_),
    .A2(_03235_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10358_ (.A1(_03218_),
    .A2(_03221_),
    .A3(_03236_),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10359_ (.A1(_03214_),
    .A2(_03237_),
    .Z(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10360_ (.A1(_03196_),
    .A2(_03238_),
    .Z(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10361_ (.A1(_03137_),
    .A2(_03151_),
    .Z(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10362_ (.A1(_03137_),
    .A2(_03151_),
    .Z(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10363_ (.A1(_03134_),
    .A2(_03240_),
    .B(_03241_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10364_ (.A1(_03139_),
    .A2(_03140_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10365_ (.A1(_03138_),
    .A2(_03141_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10366_ (.A1(_03243_),
    .A2(_03244_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10367_ (.A1(_03242_),
    .A2(_03245_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10368_ (.A1(_03082_),
    .A2(_03246_),
    .Z(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10369_ (.A1(_03239_),
    .A2(_03247_),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10370_ (.A1(_03191_),
    .A2(_03194_),
    .A3(_03248_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10371_ (.A1(_03110_),
    .A2(_03164_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10372_ (.A1(_03107_),
    .A2(_03165_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10373_ (.A1(_03250_),
    .A2(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10374_ (.A1(_03249_),
    .A2(_03252_),
    .Z(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10375_ (.I(_03169_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10376_ (.A1(_03166_),
    .A2(_03254_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10377_ (.A1(_03170_),
    .A2(_03182_),
    .B(_03255_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10378_ (.A1(_00517_),
    .A2(_03253_),
    .A3(_03256_),
    .Z(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10379_ (.A1(_03094_),
    .A2(_03184_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10380_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-4] ),
    .A2(_03183_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10381_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ),
    .A2(_03185_),
    .B1(_03183_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-4] ),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10382_ (.A1(_03259_),
    .A2(_03260_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10383_ (.A1(_03102_),
    .A2(_03258_),
    .B(_03261_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10384_ (.A1(_03257_),
    .A2(_03262_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10385_ (.A1(_03257_),
    .A2(_03262_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10386_ (.A1(_05182_),
    .A2(_03264_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10387_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[23] ),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10388_ (.A1(_05280_),
    .A2(_03266_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10389_ (.A1(_03263_),
    .A2(_03265_),
    .B(_03267_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10390_ (.A1(_03082_),
    .A2(_03246_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10391_ (.A1(_03242_),
    .A2(_03245_),
    .B(_03268_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10392_ (.A1(_03196_),
    .A2(_03238_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10393_ (.A1(_03239_),
    .A2(_03247_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10394_ (.A1(_03270_),
    .A2(_03271_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10395_ (.A1(_03198_),
    .A2(_03213_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10396_ (.A1(_03214_),
    .A2(_03237_),
    .B(_03273_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10397_ (.A1(_03200_),
    .A2(_03203_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10398_ (.A1(_03204_),
    .A2(_03212_),
    .B(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10399_ (.A1(_03037_),
    .A2(_03202_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10400_ (.A1(_03115_),
    .A2(_03277_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10401_ (.A1(net63),
    .A2(_06724_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10402_ (.A1(_02608_),
    .A2(_02704_),
    .A3(_03279_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10403_ (.A1(_03037_),
    .A2(_03280_),
    .Z(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10404_ (.A1(_03278_),
    .A2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10405_ (.A1(net63),
    .A2(_06710_),
    .B(net57),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10406_ (.A1(net63),
    .A2(_06710_),
    .A3(net57),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10407_ (.A1(_02704_),
    .A2(_03283_),
    .B(_03284_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10408_ (.A1(_00398_),
    .A2(_06708_),
    .B1(_06710_),
    .B2(_00394_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10409_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06708_),
    .A4(_06710_),
    .Z(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10410_ (.A1(_03286_),
    .A2(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10411_ (.A1(_03285_),
    .A2(_03288_),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10412_ (.A1(_03209_),
    .A2(_03289_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10413_ (.A1(_03282_),
    .A2(_03290_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10414_ (.A1(_03276_),
    .A2(_03291_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10415_ (.I(_03234_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10416_ (.A1(_03230_),
    .A2(_03293_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10417_ (.A1(_03227_),
    .A2(_03235_),
    .B(_03294_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10418_ (.A1(_03207_),
    .A2(_03210_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10419_ (.A1(_03126_),
    .A2(_03211_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10420_ (.A1(_03296_),
    .A2(_03297_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10421_ (.A1(_03232_),
    .A2(_03233_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10422_ (.A1(_03232_),
    .A2(_03233_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10423_ (.A1(_03231_),
    .A2(_03299_),
    .B(_03300_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10424_ (.A1(_00382_),
    .A2(_06742_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10425_ (.A1(_00388_),
    .A2(_06730_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10426_ (.A1(_00385_),
    .A2(_06738_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10427_ (.A1(_03302_),
    .A2(_03303_),
    .A3(_03304_),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10428_ (.A1(_03301_),
    .A2(_03305_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10429_ (.A1(_00379_),
    .A2(_00376_),
    .B(_06744_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10430_ (.A1(_00379_),
    .A2(_00376_),
    .A3(_06744_),
    .Z(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10431_ (.A1(_03307_),
    .A2(_03308_),
    .Z(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10432_ (.A1(_03138_),
    .A2(_03309_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10433_ (.I(_03310_),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10434_ (.A1(_03306_),
    .A2(_03311_),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10435_ (.A1(_03295_),
    .A2(_03298_),
    .A3(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10436_ (.A1(_03292_),
    .A2(_03313_),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10437_ (.A1(_03274_),
    .A2(_03314_),
    .Z(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10438_ (.A1(_03221_),
    .A2(_03236_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10439_ (.A1(_03221_),
    .A2(_03236_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10440_ (.A1(_03218_),
    .A2(_03316_),
    .B(_03317_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10441_ (.A1(_03138_),
    .A2(_03226_),
    .B(_03225_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10442_ (.A1(_03318_),
    .A2(_03319_),
    .Z(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10443_ (.A1(_03082_),
    .A2(_03320_),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10444_ (.A1(_03315_),
    .A2(_03321_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10445_ (.A1(_03272_),
    .A2(_03322_),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10446_ (.A1(_03269_),
    .A2(_03323_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10447_ (.A1(_03194_),
    .A2(_03248_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10448_ (.A1(_03194_),
    .A2(_03248_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10449_ (.A1(_03191_),
    .A2(_03325_),
    .B(_03326_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10450_ (.A1(_03324_),
    .A2(_03327_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10451_ (.I(_03170_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10452_ (.A1(_03329_),
    .A2(_03253_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10453_ (.A1(_03249_),
    .A2(_03252_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10454_ (.A1(_03249_),
    .A2(_03252_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10455_ (.A1(_03255_),
    .A2(_03331_),
    .B(_03332_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10456_ (.I(_03333_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10457_ (.A1(_03182_),
    .A2(_03330_),
    .B(_03334_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10458_ (.A1(_00522_),
    .A2(_03328_),
    .A3(_03335_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10459_ (.A1(_03253_),
    .A2(_03256_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10460_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-3] ),
    .A2(_03337_),
    .B(_03263_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10461_ (.A1(_03336_),
    .A2(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10462_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[24] ),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10463_ (.A1(_05280_),
    .A2(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10464_ (.A1(_05822_),
    .A2(_03339_),
    .B(_03341_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10465_ (.A1(_03094_),
    .A2(_03184_),
    .A3(_03257_),
    .A4(_03336_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10466_ (.A1(_03342_),
    .A2(_03100_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10467_ (.A1(_02681_),
    .A2(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _10468_ (.A1(_02849_),
    .A2(_02930_),
    .A3(_03096_),
    .B1(_03098_),
    .B2(_03099_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _10469_ (.A1(_03257_),
    .A2(_03336_),
    .Z(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10470_ (.A1(_03328_),
    .A2(_03335_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10471_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-3] ),
    .A2(_03337_),
    .B1(_03347_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-2] ),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10472_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-2] ),
    .A2(_03347_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _10473_ (.A1(_03259_),
    .A2(_03260_),
    .A3(_03346_),
    .B1(_03348_),
    .B2(_03349_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10474_ (.A1(_03345_),
    .A2(_03342_),
    .B(_03350_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10475_ (.A1(_03344_),
    .A2(_03351_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10476_ (.A1(_03318_),
    .A2(_03319_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10477_ (.A1(_03082_),
    .A2(_03320_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10478_ (.A1(_03353_),
    .A2(_03354_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10479_ (.A1(_03274_),
    .A2(_03314_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10480_ (.A1(_03315_),
    .A2(_03321_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10481_ (.A1(_03356_),
    .A2(_03357_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10482_ (.A1(_03276_),
    .A2(_03291_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10483_ (.A1(_03292_),
    .A2(_03313_),
    .B(_03359_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10484_ (.A1(_03278_),
    .A2(_03281_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10485_ (.A1(_03282_),
    .A2(_03290_),
    .B(_03361_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10486_ (.A1(_03037_),
    .A2(_03280_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10487_ (.A1(_03115_),
    .A2(_03363_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10488_ (.A1(net63),
    .A2(_06730_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10489_ (.A1(net57),
    .A2(_02704_),
    .A3(_03365_),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10490_ (.A1(_03037_),
    .A2(_03366_),
    .Z(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10491_ (.A1(_03364_),
    .A2(_03367_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10492_ (.A1(net63),
    .A2(_06724_),
    .B(net57),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10493_ (.A1(net63),
    .A2(_06724_),
    .A3(net57),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10494_ (.A1(_02704_),
    .A2(_03369_),
    .B(_03370_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10495_ (.A1(_00398_),
    .A2(_06710_),
    .B1(_06724_),
    .B2(_00394_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10496_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06710_),
    .A4(_06724_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10497_ (.A1(_03372_),
    .A2(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10498_ (.A1(_03371_),
    .A2(_03374_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10499_ (.A1(_03287_),
    .A2(_03375_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10500_ (.A1(_03368_),
    .A2(_03376_),
    .Z(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10501_ (.A1(_03362_),
    .A2(_03377_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10502_ (.I(_03305_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10503_ (.A1(_03301_),
    .A2(_03379_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10504_ (.A1(_03306_),
    .A2(_03311_),
    .B(_03380_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10505_ (.A1(_03285_),
    .A2(_03288_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10506_ (.A1(_03209_),
    .A2(_03289_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10507_ (.A1(_03382_),
    .A2(_03383_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10508_ (.A1(_03303_),
    .A2(_03304_),
    .Z(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10509_ (.A1(_03303_),
    .A2(_03304_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10510_ (.A1(_03302_),
    .A2(_03385_),
    .B(_03386_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10511_ (.A1(_00382_),
    .A2(_06744_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10512_ (.A1(_00388_),
    .A2(_06738_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10513_ (.A1(_00385_),
    .A2(_06742_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10514_ (.A1(_03388_),
    .A2(_03389_),
    .A3(_03390_),
    .Z(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10515_ (.A1(_03387_),
    .A2(_03391_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10516_ (.A1(_03311_),
    .A2(_03392_),
    .Z(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10517_ (.A1(_03381_),
    .A2(_03384_),
    .A3(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10518_ (.A1(_03378_),
    .A2(_03394_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10519_ (.A1(_03360_),
    .A2(_03395_),
    .Z(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10520_ (.A1(_03298_),
    .A2(_03312_),
    .Z(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10521_ (.A1(_03298_),
    .A2(_03312_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10522_ (.A1(_03295_),
    .A2(_03397_),
    .B(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10523_ (.A1(_03138_),
    .A2(_03309_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10524_ (.A1(_03308_),
    .A2(_03400_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10525_ (.A1(_03399_),
    .A2(_03401_),
    .Z(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10526_ (.A1(_03082_),
    .A2(_03402_),
    .Z(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10527_ (.A1(_03396_),
    .A2(_03403_),
    .Z(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _10528_ (.A1(_03355_),
    .A2(_03358_),
    .A3(_03404_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10529_ (.A1(_03272_),
    .A2(_03322_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10530_ (.A1(_03269_),
    .A2(_03323_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10531_ (.A1(_03406_),
    .A2(_03407_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10532_ (.I(_03408_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10533_ (.A1(_03405_),
    .A2(_03409_),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10534_ (.A1(_03324_),
    .A2(_03327_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10535_ (.A1(_03328_),
    .A2(net69),
    .B(_03411_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10536_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-1] ),
    .A2(_03410_),
    .A3(_03412_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10537_ (.A1(_03352_),
    .A2(_03413_),
    .Z(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10538_ (.A1(_03352_),
    .A2(_03413_),
    .B(_05182_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _10539_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[25] ),
    .Z(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10540_ (.A1(_05280_),
    .A2(net147),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10541_ (.A1(_03414_),
    .A2(_03415_),
    .B(_03417_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10542_ (.A1(_03399_),
    .A2(_03401_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10543_ (.A1(_03082_),
    .A2(_03402_),
    .B(_03418_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10544_ (.A1(_03360_),
    .A2(_03395_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10545_ (.A1(_03396_),
    .A2(_03403_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10546_ (.A1(_03420_),
    .A2(_03421_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10547_ (.A1(_03362_),
    .A2(_03377_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10548_ (.A1(_03378_),
    .A2(_03394_),
    .B(_03423_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10549_ (.A1(_03364_),
    .A2(_03367_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10550_ (.A1(_03368_),
    .A2(_03376_),
    .B(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10551_ (.A1(_03037_),
    .A2(_03366_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10552_ (.A1(_03115_),
    .A2(_03427_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10553_ (.A1(net63),
    .A2(_06738_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10554_ (.A1(net57),
    .A2(_02704_),
    .A3(_03429_),
    .Z(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10555_ (.A1(_03037_),
    .A2(_03430_),
    .Z(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10556_ (.A1(_03428_),
    .A2(_03431_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10557_ (.A1(net63),
    .A2(_06730_),
    .B(net57),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10558_ (.A1(net63),
    .A2(_06730_),
    .A3(net57),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10559_ (.A1(_02704_),
    .A2(_03433_),
    .B(_03434_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10560_ (.A1(_00398_),
    .A2(_06724_),
    .B1(_06730_),
    .B2(_00394_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10561_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06724_),
    .A4(_06730_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10562_ (.I(_03437_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10563_ (.A1(_03436_),
    .A2(_03438_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10564_ (.A1(_03435_),
    .A2(_03439_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10565_ (.A1(_03373_),
    .A2(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10566_ (.A1(_03432_),
    .A2(_03441_),
    .Z(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10567_ (.A1(_03426_),
    .A2(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10568_ (.I(_03391_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10569_ (.A1(_03387_),
    .A2(_03444_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10570_ (.A1(_03311_),
    .A2(_03392_),
    .B(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10571_ (.A1(_03371_),
    .A2(_03374_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10572_ (.A1(_03287_),
    .A2(_03375_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10573_ (.A1(_03447_),
    .A2(_03448_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10574_ (.A1(_03389_),
    .A2(_03390_),
    .Z(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10575_ (.A1(_03389_),
    .A2(_03390_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10576_ (.A1(_03388_),
    .A2(_03450_),
    .B(_03451_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10577_ (.A1(_00388_),
    .A2(_06742_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10578_ (.A1(_00385_),
    .A2(_06744_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10579_ (.A1(_03388_),
    .A2(_03453_),
    .A3(_03454_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10580_ (.A1(_03452_),
    .A2(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10581_ (.A1(_03311_),
    .A2(_03456_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10582_ (.A1(_03446_),
    .A2(_03449_),
    .A3(_03457_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10583_ (.A1(_03443_),
    .A2(_03458_),
    .Z(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10584_ (.A1(_03424_),
    .A2(_03459_),
    .Z(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10585_ (.A1(_03384_),
    .A2(_03393_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10586_ (.A1(_03384_),
    .A2(_03393_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10587_ (.A1(_03381_),
    .A2(_03461_),
    .B(_03462_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10588_ (.A1(_03401_),
    .A2(_03463_),
    .Z(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10589_ (.A1(_03082_),
    .A2(_03464_),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10590_ (.A1(_03460_),
    .A2(_03465_),
    .Z(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10591_ (.A1(_03422_),
    .A2(_03466_),
    .Z(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10592_ (.A1(_03419_),
    .A2(_03467_),
    .Z(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10593_ (.A1(_03358_),
    .A2(_03404_),
    .Z(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10594_ (.A1(_03358_),
    .A2(_03404_),
    .Z(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10595_ (.A1(_03355_),
    .A2(_03469_),
    .B(_03470_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10596_ (.A1(_03468_),
    .A2(_03471_),
    .Z(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10597_ (.A1(_03328_),
    .A2(_03410_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10598_ (.I(_03473_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10599_ (.A1(_03333_),
    .A2(_03473_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _10600_ (.A1(_03182_),
    .A2(_03330_),
    .A3(_03474_),
    .B(_03475_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10601_ (.A1(_03405_),
    .A2(_03409_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10602_ (.A1(_03411_),
    .A2(_03477_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10603_ (.A1(_03405_),
    .A2(_03409_),
    .B(_03478_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10604_ (.A1(_03476_),
    .A2(_03479_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10605_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ),
    .A2(_03472_),
    .A3(_03480_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10606_ (.A1(_03410_),
    .A2(_03412_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10607_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-1] ),
    .A2(_03482_),
    .B(_03414_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10608_ (.A1(_03481_),
    .A2(_03483_),
    .Z(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10609_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[26] ),
    .Z(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10610_ (.A1(_05280_),
    .A2(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10611_ (.A1(_05822_),
    .A2(_03484_),
    .B(_03486_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10612_ (.A1(_03422_),
    .A2(_03466_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10613_ (.I(_03419_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10614_ (.A1(_03488_),
    .A2(_03467_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10615_ (.A1(_03082_),
    .A2(_03464_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10616_ (.A1(_03401_),
    .A2(_03463_),
    .B(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10617_ (.A1(_03424_),
    .A2(_03459_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10618_ (.A1(_03460_),
    .A2(_03465_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10619_ (.A1(_03492_),
    .A2(_03493_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10620_ (.A1(_03426_),
    .A2(_03442_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10621_ (.A1(_03443_),
    .A2(_03458_),
    .B(_03495_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10622_ (.A1(_03428_),
    .A2(_03431_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10623_ (.A1(_03432_),
    .A2(_03441_),
    .B(_03497_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10624_ (.A1(net63),
    .A2(_06738_),
    .B(net57),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10625_ (.A1(net63),
    .A2(_06738_),
    .A3(net57),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10626_ (.A1(_02704_),
    .A2(_03499_),
    .B(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10627_ (.A1(_00398_),
    .A2(_06730_),
    .B1(_06738_),
    .B2(_00394_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10628_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06730_),
    .A4(_06738_),
    .Z(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10629_ (.A1(_03502_),
    .A2(_03503_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10630_ (.A1(_03437_),
    .A2(_03501_),
    .A3(_03504_),
    .Z(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10631_ (.A1(_03037_),
    .A2(_03430_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10632_ (.A1(_03115_),
    .A2(_03506_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10633_ (.A1(net63),
    .A2(_06742_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10634_ (.A1(net57),
    .A2(_02704_),
    .A3(_03508_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10635_ (.A1(_03037_),
    .A2(_03509_),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10636_ (.A1(_03507_),
    .A2(_03510_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10637_ (.A1(_03505_),
    .A2(_03511_),
    .Z(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10638_ (.A1(_03498_),
    .A2(_03512_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10639_ (.A1(_03452_),
    .A2(_03455_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10640_ (.A1(_03311_),
    .A2(_03456_),
    .B(_03514_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10641_ (.A1(_03435_),
    .A2(_03439_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10642_ (.A1(_03373_),
    .A2(_03440_),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10643_ (.A1(_03516_),
    .A2(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10644_ (.A1(_00388_),
    .A2(_00385_),
    .B(_06744_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10645_ (.A1(_00388_),
    .A2(_00385_),
    .A3(_06744_),
    .Z(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10646_ (.A1(_03519_),
    .A2(_03520_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10647_ (.A1(_03453_),
    .A2(_03454_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10648_ (.A1(_03453_),
    .A2(_03454_),
    .Z(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10649_ (.A1(_00382_),
    .A2(_03522_),
    .B1(_03523_),
    .B2(_03388_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10650_ (.A1(_03521_),
    .A2(_03524_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10651_ (.A1(_03311_),
    .A2(_03525_),
    .Z(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10652_ (.A1(_03515_),
    .A2(_03518_),
    .A3(_03526_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10653_ (.A1(_03513_),
    .A2(_03527_),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10654_ (.A1(_03496_),
    .A2(_03528_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10655_ (.A1(_03449_),
    .A2(_03457_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10656_ (.A1(_03449_),
    .A2(_03457_),
    .Z(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10657_ (.A1(_03446_),
    .A2(_03530_),
    .B(_03531_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10658_ (.A1(_03401_),
    .A2(_03532_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10659_ (.A1(_03082_),
    .A2(_03533_),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10660_ (.A1(_03529_),
    .A2(_03534_),
    .Z(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10661_ (.A1(_03494_),
    .A2(_03535_),
    .Z(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10662_ (.A1(_03491_),
    .A2(_03536_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10663_ (.A1(_03487_),
    .A2(_03489_),
    .B(_03537_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10664_ (.A1(_03487_),
    .A2(_03489_),
    .A3(_03537_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10665_ (.A1(_03538_),
    .A2(_03539_),
    .Z(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10666_ (.A1(_03468_),
    .A2(_03471_),
    .Z(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10667_ (.A1(_03476_),
    .A2(_03479_),
    .B(_03472_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10668_ (.A1(_03541_),
    .A2(_03542_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10669_ (.A1(_00537_),
    .A2(_03540_),
    .A3(_03543_),
    .Z(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10670_ (.A1(_03345_),
    .A2(net79),
    .B1(_03343_),
    .B2(_02681_),
    .C(_03350_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10671_ (.A1(_03413_),
    .A2(_03481_),
    .Z(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10672_ (.I(_03546_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10673_ (.A1(_03472_),
    .A2(_03480_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10674_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ),
    .A2(_03548_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10675_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-1] ),
    .A2(_03482_),
    .B1(_03548_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10676_ (.A1(_03549_),
    .A2(_03550_),
    .Z(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10677_ (.A1(_03545_),
    .A2(_03547_),
    .B(_03551_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10678_ (.A1(_03544_),
    .A2(_03552_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10679_ (.A1(_03544_),
    .A2(_03552_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10680_ (.A1(_05182_),
    .A2(_03554_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10681_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[27] ),
    .Z(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10682_ (.A1(_05280_),
    .A2(_03556_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10683_ (.A1(_03553_),
    .A2(_03555_),
    .B(_03557_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10684_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[28] ),
    .Z(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10685_ (.A1(_03082_),
    .A2(_03533_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10686_ (.A1(_03401_),
    .A2(_03532_),
    .B(_03559_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10687_ (.A1(_03496_),
    .A2(_03528_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10688_ (.A1(_03529_),
    .A2(_03534_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10689_ (.A1(_03561_),
    .A2(_03562_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10690_ (.A1(_03498_),
    .A2(_03512_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10691_ (.A1(_03513_),
    .A2(_03527_),
    .B(_03564_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10692_ (.A1(_03507_),
    .A2(_03510_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10693_ (.A1(_03505_),
    .A2(_03511_),
    .B(_03566_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10694_ (.A1(net63),
    .A2(_06742_),
    .B(net57),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10695_ (.A1(net63),
    .A2(_06742_),
    .A3(net57),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10696_ (.A1(_02704_),
    .A2(_03568_),
    .B(_03569_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10697_ (.A1(_00398_),
    .A2(_06738_),
    .B1(_06742_),
    .B2(_00394_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10698_ (.A1(_00398_),
    .A2(_00394_),
    .A3(_06738_),
    .A4(_06742_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10699_ (.A1(_03571_),
    .A2(_03572_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10700_ (.A1(_03570_),
    .A2(_03573_),
    .Z(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10701_ (.A1(_03503_),
    .A2(_03574_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10702_ (.A1(_03037_),
    .A2(_03509_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10703_ (.A1(_03115_),
    .A2(_03576_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10704_ (.A1(net63),
    .A2(_06744_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10705_ (.A1(net57),
    .A2(_02704_),
    .A3(_03578_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10706_ (.A1(_03037_),
    .A2(_03579_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10707_ (.A1(_03577_),
    .A2(_03580_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10708_ (.I(_03581_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10709_ (.A1(_03575_),
    .A2(_03582_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10710_ (.A1(_03567_),
    .A2(_03583_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10711_ (.A1(_00382_),
    .A2(_03520_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10712_ (.A1(_03311_),
    .A2(_03525_),
    .B(_03585_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10713_ (.A1(_03501_),
    .A2(_03504_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10714_ (.A1(_03501_),
    .A2(_03504_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10715_ (.A1(_03437_),
    .A2(_03587_),
    .B(_03588_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10716_ (.A1(_03388_),
    .A2(_03519_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10717_ (.A1(_03585_),
    .A2(_03590_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10718_ (.A1(_03311_),
    .A2(_03591_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10719_ (.A1(_03589_),
    .A2(_03592_),
    .Z(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10720_ (.A1(_03586_),
    .A2(_03593_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10721_ (.A1(_03584_),
    .A2(_03594_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10722_ (.A1(_03565_),
    .A2(_03595_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10723_ (.A1(_03518_),
    .A2(_03526_),
    .Z(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10724_ (.A1(_03518_),
    .A2(_03526_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10725_ (.A1(_03515_),
    .A2(_03597_),
    .B(_03598_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10726_ (.A1(_03401_),
    .A2(_03599_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10727_ (.A1(_03082_),
    .A2(_03600_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10728_ (.A1(_03596_),
    .A2(_03601_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10729_ (.I(_03602_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10730_ (.A1(_03563_),
    .A2(_03603_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10731_ (.A1(_03560_),
    .A2(_03604_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10732_ (.A1(_03494_),
    .A2(_03535_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10733_ (.A1(_03491_),
    .A2(_03536_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10734_ (.A1(_03606_),
    .A2(_03607_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10735_ (.A1(_03605_),
    .A2(_03608_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10736_ (.I(_03541_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10737_ (.I(_03539_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10738_ (.A1(_03610_),
    .A2(_03538_),
    .B(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10739_ (.I(_03540_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10740_ (.A1(_03476_),
    .A2(_03479_),
    .B(_03613_),
    .C(_03472_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10741_ (.A1(_03612_),
    .A2(_03614_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _10742_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[2] ),
    .A2(_03609_),
    .A3(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10743_ (.A1(_03613_),
    .A2(_03543_),
    .Z(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10744_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[1] ),
    .A2(_03617_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10745_ (.A1(_03618_),
    .A2(_03554_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10746_ (.A1(_03616_),
    .A2(_03619_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10747_ (.I0(_03558_),
    .I1(_03620_),
    .S(_05171_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10748_ (.I(_03621_),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10749_ (.A1(_03544_),
    .A2(_03616_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10750_ (.A1(_03609_),
    .A2(_03615_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10751_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[1] ),
    .A2(_03617_),
    .B1(_03623_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[2] ),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10752_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[2] ),
    .A2(_03623_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10753_ (.A1(_03544_),
    .A2(_03546_),
    .A3(_03616_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _10754_ (.A1(_03551_),
    .A2(_03622_),
    .B1(_03624_),
    .B2(_03625_),
    .C1(_03626_),
    .C2(_03545_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10755_ (.A1(_03082_),
    .A2(_03600_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10756_ (.A1(_03401_),
    .A2(_03599_),
    .B(_03628_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10757_ (.A1(_03565_),
    .A2(_03595_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10758_ (.A1(_03596_),
    .A2(_03601_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10759_ (.A1(_03630_),
    .A2(_03631_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10760_ (.A1(_03567_),
    .A2(_03583_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10761_ (.A1(_03584_),
    .A2(_03594_),
    .B(_03633_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10762_ (.A1(_03577_),
    .A2(_03580_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10763_ (.A1(_03575_),
    .A2(_03582_),
    .B(_03635_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10764_ (.A1(_03037_),
    .A2(_03579_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10765_ (.A1(_03031_),
    .A2(_03579_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10766_ (.A1(_03031_),
    .A2(_03637_),
    .B(_03638_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10767_ (.A1(net58),
    .A2(net63),
    .B(_06744_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10768_ (.A1(net58),
    .A2(net63),
    .A3(_06744_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10769_ (.A1(_02704_),
    .A2(_03640_),
    .B(_03641_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10770_ (.A1(_00398_),
    .A2(_06742_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10771_ (.A1(_00394_),
    .A2(_06744_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10772_ (.A1(_03643_),
    .A2(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10773_ (.I(_03644_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10774_ (.A1(_00398_),
    .A2(_06742_),
    .A3(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10775_ (.A1(_03645_),
    .A2(_03647_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10776_ (.A1(_03642_),
    .A2(_03648_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10777_ (.A1(_03572_),
    .A2(_03649_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10778_ (.A1(_03639_),
    .A2(_03650_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10779_ (.A1(_03636_),
    .A2(_03651_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10780_ (.A1(_03388_),
    .A2(_03519_),
    .Z(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10781_ (.A1(_03311_),
    .A2(_03653_),
    .B(_03585_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10782_ (.A1(_03570_),
    .A2(_03573_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10783_ (.A1(_03503_),
    .A2(_03574_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10784_ (.A1(_03655_),
    .A2(_03656_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10785_ (.A1(_03592_),
    .A2(_03657_),
    .Z(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10786_ (.A1(_03654_),
    .A2(_03658_),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10787_ (.A1(_03652_),
    .A2(_03659_),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10788_ (.A1(_03634_),
    .A2(_03660_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10789_ (.A1(_03589_),
    .A2(_03592_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10790_ (.A1(_03586_),
    .A2(_03593_),
    .B(_03662_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10791_ (.A1(_03401_),
    .A2(_03663_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10792_ (.A1(_03082_),
    .A2(_03664_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10793_ (.A1(_03661_),
    .A2(_03665_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10794_ (.A1(_03629_),
    .A2(_03632_),
    .A3(_03666_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10795_ (.A1(_03563_),
    .A2(_03603_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10796_ (.A1(_03560_),
    .A2(_03604_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10797_ (.A1(_03668_),
    .A2(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10798_ (.A1(_03606_),
    .A2(_03607_),
    .B(_03605_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10799_ (.A1(_03612_),
    .A2(_03614_),
    .B(_03609_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10800_ (.A1(_03671_),
    .A2(_03672_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _10801_ (.A1(_03667_),
    .A2(_03670_),
    .A3(_03673_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10802_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[3] ),
    .A2(_03674_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10803_ (.A1(_03627_),
    .A2(_03675_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10804_ (.A1(_03627_),
    .A2(_03675_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10805_ (.A1(_05182_),
    .A2(_03677_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10806_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[29] ),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10807_ (.A1(_05280_),
    .A2(_03679_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10808_ (.A1(_03676_),
    .A2(_03678_),
    .B(_03680_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10809_ (.A1(_03668_),
    .A2(_03669_),
    .B(_03667_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10810_ (.A1(_03668_),
    .A2(_03669_),
    .A3(_03667_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10811_ (.A1(_03681_),
    .A2(_03673_),
    .B(_03682_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10812_ (.A1(_03632_),
    .A2(_03666_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10813_ (.A1(_03632_),
    .A2(_03666_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10814_ (.A1(_03629_),
    .A2(_03684_),
    .B(_03685_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10815_ (.A1(_03082_),
    .A2(_03664_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10816_ (.A1(_03401_),
    .A2(_03663_),
    .B(_03687_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10817_ (.A1(_03634_),
    .A2(_03660_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10818_ (.A1(_03661_),
    .A2(_03665_),
    .B(_03689_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10819_ (.A1(_03592_),
    .A2(_03657_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10820_ (.A1(_03654_),
    .A2(_03658_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10821_ (.A1(_03691_),
    .A2(_03692_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10822_ (.I(_03693_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10823_ (.A1(_03401_),
    .A2(_03694_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10824_ (.A1(_03082_),
    .A2(_03695_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10825_ (.A1(_03636_),
    .A2(_03651_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10826_ (.A1(_03652_),
    .A2(_03659_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10827_ (.A1(_03697_),
    .A2(_03698_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10828_ (.A1(_03642_),
    .A2(_03645_),
    .A3(_03647_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10829_ (.A1(_03572_),
    .A2(_03649_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10830_ (.A1(_03700_),
    .A2(_03701_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10831_ (.A1(_03592_),
    .A2(_03702_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10832_ (.A1(_03654_),
    .A2(_03703_),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10833_ (.A1(_03639_),
    .A2(_03650_),
    .B(_03638_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10834_ (.I(_03705_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10835_ (.A1(_00398_),
    .A2(_00394_),
    .B(_06744_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10836_ (.A1(_00398_),
    .A2(_03646_),
    .B(_03707_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10837_ (.A1(_03642_),
    .A2(_03708_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10838_ (.A1(_03647_),
    .A2(_03709_),
    .Z(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10839_ (.A1(_03639_),
    .A2(_03710_),
    .Z(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10840_ (.A1(_03706_),
    .A2(_03711_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10841_ (.A1(_03704_),
    .A2(_03712_),
    .Z(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10842_ (.A1(_03699_),
    .A2(_03713_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10843_ (.A1(_03696_),
    .A2(_03714_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10844_ (.A1(_03688_),
    .A2(_03690_),
    .A3(_03715_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10845_ (.A1(_03686_),
    .A2(_03716_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10846_ (.A1(_03686_),
    .A2(_03716_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10847_ (.A1(_03717_),
    .A2(_03718_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10848_ (.A1(_03683_),
    .A2(_03719_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10849_ (.A1(_00552_),
    .A2(_03720_),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10850_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[3] ),
    .A2(_03674_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10851_ (.A1(_03722_),
    .A2(_03677_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10852_ (.A1(_03721_),
    .A2(_03723_),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10853_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[30] ),
    .Z(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10854_ (.A1(_05280_),
    .A2(_03725_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10855_ (.A1(_05822_),
    .A2(_03724_),
    .B(_03726_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10856_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[31] ),
    .Z(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10857_ (.A1(_03683_),
    .A2(_03719_),
    .B(_03717_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10858_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[5] ),
    .A2(_03728_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10859_ (.A1(_03592_),
    .A2(_03702_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10860_ (.A1(_03654_),
    .A2(_03703_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10861_ (.A1(_03730_),
    .A2(_03731_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10862_ (.A1(_03401_),
    .A2(_03707_),
    .A3(_03732_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10863_ (.A1(_03690_),
    .A2(_03715_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10864_ (.A1(_03690_),
    .A2(_03715_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10865_ (.A1(_03688_),
    .A2(_03734_),
    .B(_03735_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10866_ (.A1(_03704_),
    .A2(_03712_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10867_ (.A1(_03706_),
    .A2(_03711_),
    .B(_03737_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10868_ (.A1(_03699_),
    .A2(_03713_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10869_ (.A1(_03696_),
    .A2(_03714_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10870_ (.A1(_03739_),
    .A2(_03740_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10871_ (.A1(_03642_),
    .A2(_03708_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10872_ (.A1(_03647_),
    .A2(_03709_),
    .B(_03742_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10873_ (.A1(_03082_),
    .A2(_03695_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10874_ (.A1(_03401_),
    .A2(_03694_),
    .B(_03744_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10875_ (.A1(_03031_),
    .A2(_03637_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10876_ (.A1(_03746_),
    .A2(_03710_),
    .B(_03638_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10877_ (.A1(_03311_),
    .A2(_03585_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10878_ (.A1(_03311_),
    .A2(_03653_),
    .B(_03748_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10879_ (.A1(_03747_),
    .A2(_03749_),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10880_ (.A1(_03743_),
    .A2(_03745_),
    .A3(_03750_),
    .Z(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10881_ (.A1(_03082_),
    .A2(_03741_),
    .A3(_03751_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10882_ (.A1(_03736_),
    .A2(_03738_),
    .A3(_03752_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10883_ (.A1(_03642_),
    .A2(_03733_),
    .A3(_03753_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10884_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[3] ),
    .A2(_03674_),
    .B1(_03720_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[4] ),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10885_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[4] ),
    .A2(_03720_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10886_ (.A1(_03677_),
    .A2(_03721_),
    .B1(_03755_),
    .B2(_03756_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10887_ (.A1(_03729_),
    .A2(_03754_),
    .A3(_03757_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10888_ (.I0(_03727_),
    .I1(_03758_),
    .S(_05171_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10889_ (.I(_03759_),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10890_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-25] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-25] ),
    .S(_05171_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10891_ (.I(_03760_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10892_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-24] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-24] ),
    .S(_05171_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10893_ (.I(_03761_),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10894_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-23] ),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10895_ (.A1(_05822_),
    .A2(_06765_),
    .B(_03762_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10896_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-22] ),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10897_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-22] ),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10898_ (.A1(_05387_),
    .A2(_03763_),
    .B(_03764_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10899_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-21] ),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10900_ (.A1(_05822_),
    .A2(_06777_),
    .B(_03765_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10901_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-20] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-20] ),
    .S(_05171_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10902_ (.I(_03766_),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10903_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-19] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-19] ),
    .S(_05171_),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10904_ (.I(_03767_),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10905_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-18] ),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10906_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-18] ),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10907_ (.A1(_05387_),
    .A2(_03768_),
    .B(_03769_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10908_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-17] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-17] ),
    .S(_05171_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10909_ (.I(_03770_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10910_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-16] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-16] ),
    .S(_05171_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10911_ (.I(_03771_),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10912_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-15] ),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10913_ (.A1(_05822_),
    .A2(_06811_),
    .B(_03772_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10914_ (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-14] ),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10915_ (.A1(_05387_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-14] ),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10916_ (.A1(_05387_),
    .A2(_03773_),
    .B(_03774_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10917_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-13] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-13] ),
    .S(_05171_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10918_ (.I(_03775_),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10919_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-12] ),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10920_ (.A1(_05822_),
    .A2(_06824_),
    .B(_03776_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10921_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-11] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-11] ),
    .S(_05171_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10922_ (.I(_03777_),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10923_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-10] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-10] ),
    .S(_05171_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10924_ (.I(_03778_),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10925_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-9] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-9] ),
    .S(_05171_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10926_ (.I(_03779_),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10927_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-8] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-8] ),
    .S(_05171_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10928_ (.I(_03780_),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10929_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-7] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-7] ),
    .S(_05171_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10930_ (.I(_03781_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10931_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-6] ),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10932_ (.A1(_05822_),
    .A2(_00312_),
    .B(_03782_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10933_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-5] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-5] ),
    .S(_05171_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10934_ (.I(_03783_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10935_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-4] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-4] ),
    .S(_05171_),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10936_ (.I(_03784_),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10937_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-3] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-3] ),
    .S(_05171_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10938_ (.I(_03785_),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10939_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-2] ),
    .S(_05171_),
    .Z(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10940_ (.I(_03786_),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10941_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-1] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-1] ),
    .S(_05171_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10942_ (.I(_03787_),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10943_ (.I0(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[0] ),
    .I1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[0] ),
    .S(_05171_),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10944_ (.I(_03788_),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10945_ (.A1(_05280_),
    .A2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[1] ),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10946_ (.A1(_05822_),
    .A2(_00346_),
    .B(_03789_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10947_ (.A1(_00390_),
    .A2(_02409_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10948_ (.A1(_00393_),
    .A2(_02238_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10949_ (.A1(_03790_),
    .A2(_03791_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10950_ (.A1(_03790_),
    .A2(_03791_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10951_ (.A1(_00397_),
    .A2(_02236_),
    .A3(_03793_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10952_ (.A1(_00387_),
    .A2(_02238_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10953_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02499_),
    .A4(_02409_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10954_ (.A1(_00381_),
    .A2(_02499_),
    .B1(_02409_),
    .B2(_00384_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10955_ (.A1(_03796_),
    .A2(_03797_),
    .Z(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10956_ (.I(_03796_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10957_ (.A1(_03795_),
    .A2(_03798_),
    .B(_03799_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10958_ (.A1(_00387_),
    .A2(_02409_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10959_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02584_),
    .A4(_02499_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10960_ (.A1(_00381_),
    .A2(net135),
    .B1(_02499_),
    .B2(_00384_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10961_ (.A1(_03802_),
    .A2(_03803_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10962_ (.A1(_03801_),
    .A2(_03804_),
    .Z(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10963_ (.A1(_03800_),
    .A2(_03805_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10964_ (.A1(_00397_),
    .A2(_02153_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10965_ (.A1(_00390_),
    .A2(_02238_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10966_ (.A1(_00393_),
    .A2(_02236_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10967_ (.A1(_03808_),
    .A2(_03809_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10968_ (.A1(_03807_),
    .A2(_03810_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10969_ (.A1(_03795_),
    .A2(_03798_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10970_ (.A1(_03796_),
    .A2(_03812_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10971_ (.A1(_03813_),
    .A2(_03805_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10972_ (.A1(_03806_),
    .A2(_03811_),
    .B(_03814_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10973_ (.A1(_00378_),
    .A2(net135),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10974_ (.I(_03816_),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10975_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02762_),
    .A4(_02586_),
    .Z(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10976_ (.A1(_00372_),
    .A2(_02762_),
    .B1(_02586_),
    .B2(_00375_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10977_ (.A1(_03818_),
    .A2(_03819_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10978_ (.A1(_03817_),
    .A2(_03820_),
    .B(_03818_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10979_ (.A1(_00361_),
    .A2(_02940_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10980_ (.A1(_00365_),
    .A2(_02938_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10981_ (.A1(_03822_),
    .A2(_03823_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10982_ (.A1(_00369_),
    .A2(_02854_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10983_ (.A1(_03822_),
    .A2(_03823_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10984_ (.A1(_03824_),
    .A2(_03825_),
    .B(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10985_ (.A1(_00378_),
    .A2(_02586_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10986_ (.I(_03828_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10987_ (.A1(_00372_),
    .A2(_02854_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10988_ (.A1(_00375_),
    .A2(_02762_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10989_ (.A1(_03829_),
    .A2(_03830_),
    .A3(_03831_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10990_ (.A1(_03827_),
    .A2(_03832_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10991_ (.A1(_03827_),
    .A2(_03832_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10992_ (.A1(_03821_),
    .A2(_03833_),
    .B(_03834_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10993_ (.A1(_03802_),
    .A2(_03801_),
    .A3(_03803_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10994_ (.A1(_03802_),
    .A2(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10995_ (.A1(_00387_),
    .A2(_02499_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10996_ (.A1(_00381_),
    .A2(_02586_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10997_ (.A1(_00384_),
    .A2(net135),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10998_ (.A1(_03838_),
    .A2(_03839_),
    .A3(_03840_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10999_ (.A1(_03837_),
    .A2(_03841_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11000_ (.A1(_00397_),
    .A2(_02236_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11001_ (.A1(_03843_),
    .A2(_03793_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11002_ (.A1(_03842_),
    .A2(_03844_),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11003_ (.A1(_03835_),
    .A2(_03845_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11004_ (.A1(_03835_),
    .A2(_03845_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11005_ (.A1(_03815_),
    .A2(_03846_),
    .B(_03847_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11006_ (.A1(_03792_),
    .A2(_03794_),
    .B(_03848_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11007_ (.I(_03849_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11008_ (.A1(_03792_),
    .A2(_03794_),
    .A3(_03848_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11009_ (.A1(_03849_),
    .A2(_03851_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11010_ (.A1(_03835_),
    .A2(_03845_),
    .A3(_03815_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11011_ (.A1(_03821_),
    .A2(_03833_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11012_ (.A1(_00359_),
    .A2(_02940_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11013_ (.A1(net66),
    .A2(_03189_),
    .B1(_03018_),
    .B2(net83),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11014_ (.A1(net66),
    .A2(net83),
    .A3(_03189_),
    .A4(_03018_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11015_ (.A1(_03855_),
    .A2(_03856_),
    .B(_03857_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11016_ (.A1(_00359_),
    .A2(_03018_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11017_ (.A1(_00351_),
    .A2(_03266_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11018_ (.A1(net83),
    .A2(_03189_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11019_ (.A1(_03859_),
    .A2(_03860_),
    .A3(_03861_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11020_ (.A1(_03858_),
    .A2(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11021_ (.A1(_03822_),
    .A2(_03823_),
    .A3(_03825_),
    .Z(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11022_ (.A1(_03858_),
    .A2(_03862_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11023_ (.A1(_03863_),
    .A2(_03864_),
    .B(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11024_ (.A1(_00369_),
    .A2(_02938_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11025_ (.A1(_00365_),
    .A2(_02940_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11026_ (.A1(_00361_),
    .A2(_03018_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11027_ (.A1(_03867_),
    .A2(_03868_),
    .A3(_03869_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11028_ (.A1(net66),
    .A2(_03266_),
    .B1(_03189_),
    .B2(net54),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11029_ (.A1(net66),
    .A2(net54),
    .A3(_03266_),
    .A4(_03189_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11030_ (.A1(_03859_),
    .A2(_03871_),
    .B(_03872_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11031_ (.A1(_00359_),
    .A2(_03189_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11032_ (.A1(net87),
    .A2(_03340_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11033_ (.A1(net83),
    .A2(_03266_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11034_ (.A1(_03874_),
    .A2(_03875_),
    .A3(_03876_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11035_ (.A1(_03877_),
    .A2(_03873_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11036_ (.A1(_03870_),
    .A2(_03878_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11037_ (.A1(_03866_),
    .A2(_03879_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11038_ (.A1(_03866_),
    .A2(_03879_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11039_ (.A1(_03854_),
    .A2(_03880_),
    .B(_03881_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11040_ (.A1(_03830_),
    .A2(_03831_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11041_ (.A1(_03830_),
    .A2(_03831_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11042_ (.A1(_03829_),
    .A2(_03883_),
    .B(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11043_ (.A1(_03868_),
    .A2(_03869_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11044_ (.A1(_03868_),
    .A2(_03869_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11045_ (.A1(_03867_),
    .A2(_03886_),
    .B(_03887_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11046_ (.A1(_00378_),
    .A2(_02762_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11047_ (.I(_03889_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11048_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02938_),
    .A4(_02854_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11049_ (.A1(_00372_),
    .A2(_02938_),
    .B1(_02854_),
    .B2(_00375_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11050_ (.A1(_03891_),
    .A2(_03892_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11051_ (.A1(_03890_),
    .A2(_03893_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11052_ (.A1(_03888_),
    .A2(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11053_ (.A1(_03885_),
    .A2(_03895_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11054_ (.A1(_03873_),
    .A2(_03877_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11055_ (.A1(_03870_),
    .A2(_03878_),
    .B(_03897_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11056_ (.A1(_00369_),
    .A2(_02940_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11057_ (.A1(_00361_),
    .A2(_03189_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11058_ (.A1(_00365_),
    .A2(_03018_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11059_ (.A1(_03899_),
    .A2(_03900_),
    .A3(_03901_),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11060_ (.A1(net66),
    .A2(_03340_),
    .B1(_03266_),
    .B2(net54),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11061_ (.A1(net66),
    .A2(net54),
    .A3(_03340_),
    .A4(_03266_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11062_ (.A1(_03874_),
    .A2(_03903_),
    .B(_03904_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11063_ (.A1(_00359_),
    .A2(_03266_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11064_ (.A1(net87),
    .A2(_03416_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11065_ (.A1(net54),
    .A2(_03340_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11066_ (.A1(_03906_),
    .A2(_03907_),
    .A3(_03908_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11067_ (.A1(_03905_),
    .A2(_03909_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11068_ (.A1(_03902_),
    .A2(_03910_),
    .Z(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11069_ (.A1(_03896_),
    .A2(_03898_),
    .A3(_03911_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11070_ (.A1(_03882_),
    .A2(_03912_),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11071_ (.A1(_03882_),
    .A2(_03912_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11072_ (.A1(_03853_),
    .A2(_03913_),
    .B(_03914_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11073_ (.A1(_03898_),
    .A2(_03911_),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11074_ (.A1(_03898_),
    .A2(_03911_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11075_ (.A1(_03896_),
    .A2(_03916_),
    .B(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11076_ (.A1(_03890_),
    .A2(_03893_),
    .B(_03891_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11077_ (.A1(_03900_),
    .A2(_03901_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11078_ (.A1(_03900_),
    .A2(_03901_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11079_ (.A1(_03899_),
    .A2(_03920_),
    .B(_03921_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11080_ (.A1(_00378_),
    .A2(_02854_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11081_ (.I(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11082_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02940_),
    .A4(_02938_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11083_ (.A1(_00372_),
    .A2(_02940_),
    .B1(_02938_),
    .B2(_00375_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11084_ (.A1(_03925_),
    .A2(_03926_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11085_ (.A1(_03924_),
    .A2(_03927_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11086_ (.A1(_03922_),
    .A2(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11087_ (.A1(_03919_),
    .A2(_03929_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11088_ (.A1(_03905_),
    .A2(_03909_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11089_ (.A1(_03902_),
    .A2(_03910_),
    .B(_03931_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11090_ (.A1(_00369_),
    .A2(_03018_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11091_ (.A1(_00361_),
    .A2(_03266_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11092_ (.A1(_00365_),
    .A2(_03189_),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11093_ (.A1(_03933_),
    .A2(_03934_),
    .A3(_03935_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11094_ (.A1(net86),
    .A2(_03416_),
    .B1(_03340_),
    .B2(net83),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11095_ (.A1(net86),
    .A2(net83),
    .A3(_03416_),
    .A4(_03340_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11096_ (.A1(_03906_),
    .A2(_03937_),
    .B(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11097_ (.A1(_00359_),
    .A2(_03340_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11098_ (.A1(_00351_),
    .A2(_03485_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11099_ (.A1(net84),
    .A2(_03416_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11100_ (.A1(_03940_),
    .A2(_03941_),
    .A3(_03942_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11101_ (.A1(_03939_),
    .A2(_03943_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11102_ (.A1(_03936_),
    .A2(_03944_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11103_ (.A1(_03932_),
    .A2(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11104_ (.A1(_03930_),
    .A2(_03946_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11105_ (.A1(_03918_),
    .A2(_03947_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11106_ (.A1(_03842_),
    .A2(_03844_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11107_ (.A1(_03837_),
    .A2(_03841_),
    .B(_03949_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11108_ (.A1(_03888_),
    .A2(_03894_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11109_ (.A1(_03885_),
    .A2(_03895_),
    .B(_03951_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11110_ (.A1(_03839_),
    .A2(_03840_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11111_ (.A1(_03839_),
    .A2(_03840_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11112_ (.A1(_03838_),
    .A2(_03953_),
    .B(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11113_ (.A1(_00387_),
    .A2(net135),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11114_ (.A1(_00384_),
    .A2(_02586_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11115_ (.A1(_02762_),
    .A2(_00381_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11116_ (.A1(_03956_),
    .A2(_03957_),
    .A3(_03958_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11117_ (.A1(_03955_),
    .A2(_03959_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11118_ (.A1(_00397_),
    .A2(_02238_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11119_ (.A1(_00393_),
    .A2(_02409_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11120_ (.A1(_00390_),
    .A2(_02499_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11121_ (.A1(_03962_),
    .A2(_03963_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11122_ (.A1(_03961_),
    .A2(_03964_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11123_ (.A1(_03960_),
    .A2(_03965_),
    .Z(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11124_ (.A1(_03950_),
    .A2(_03952_),
    .A3(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11125_ (.A1(_03948_),
    .A2(_03967_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11126_ (.A1(_03915_),
    .A2(_03968_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11127_ (.A1(_03915_),
    .A2(_03968_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11128_ (.A1(_03852_),
    .A2(_03969_),
    .B(_03970_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11129_ (.A1(_03962_),
    .A2(_03963_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11130_ (.A1(_00397_),
    .A2(_02238_),
    .A3(_03964_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11131_ (.A1(_03952_),
    .A2(_03966_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11132_ (.A1(_03952_),
    .A2(_03966_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11133_ (.A1(_03950_),
    .A2(_03974_),
    .B(_03975_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11134_ (.A1(_03972_),
    .A2(_03973_),
    .B(_03976_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11135_ (.A1(_03972_),
    .A2(_03973_),
    .A3(_03976_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11136_ (.A1(_03977_),
    .A2(_03978_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11137_ (.A1(_03918_),
    .A2(_03947_),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11138_ (.A1(_03948_),
    .A2(_03967_),
    .B(_03980_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11139_ (.A1(_03932_),
    .A2(_03945_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11140_ (.A1(_03930_),
    .A2(_03946_),
    .B(_03982_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11141_ (.A1(_03939_),
    .A2(_03943_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11142_ (.A1(_03936_),
    .A2(_03944_),
    .B(_03984_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11143_ (.A1(net86),
    .A2(_03485_),
    .B1(_03416_),
    .B2(net84),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11144_ (.A1(net86),
    .A2(net84),
    .A3(_03485_),
    .A4(_03416_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11145_ (.A1(_03940_),
    .A2(_03986_),
    .B(_03987_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11146_ (.A1(_00359_),
    .A2(_03416_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11147_ (.A1(_03556_),
    .A2(_00351_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11148_ (.A1(net84),
    .A2(_03485_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11149_ (.A1(_03989_),
    .A2(_03990_),
    .A3(_03991_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11150_ (.A1(_03988_),
    .A2(_03992_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11151_ (.A1(_00369_),
    .A2(_03189_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11152_ (.A1(_03340_),
    .A2(_00361_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11153_ (.A1(_00365_),
    .A2(_03266_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11154_ (.A1(_03994_),
    .A2(_03995_),
    .A3(_03996_),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11155_ (.A1(_03997_),
    .A2(_03993_),
    .Z(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11156_ (.A1(_03985_),
    .A2(_03998_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11157_ (.A1(_03924_),
    .A2(_03927_),
    .B(_03925_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11158_ (.A1(_03934_),
    .A2(_03935_),
    .Z(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11159_ (.A1(_03934_),
    .A2(_03935_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11160_ (.A1(_03933_),
    .A2(_04001_),
    .B(_04002_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11161_ (.A1(_00378_),
    .A2(_02938_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11162_ (.I(_04004_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11163_ (.A1(_00375_),
    .A2(_02940_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11164_ (.A1(_03018_),
    .A2(_00372_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11165_ (.A1(_04005_),
    .A2(_04006_),
    .A3(_04007_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11166_ (.A1(_04003_),
    .A2(_04008_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11167_ (.A1(_04000_),
    .A2(_04009_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11168_ (.A1(_03999_),
    .A2(_04010_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11169_ (.A1(_03983_),
    .A2(_04011_),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11170_ (.I(_03959_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11171_ (.A1(_03955_),
    .A2(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11172_ (.A1(_03960_),
    .A2(_03965_),
    .B(_04014_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11173_ (.A1(_03922_),
    .A2(_03928_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11174_ (.A1(_03919_),
    .A2(_03929_),
    .B(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11175_ (.A1(_00397_),
    .A2(_02409_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11176_ (.A1(_00393_),
    .A2(_02499_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11177_ (.A1(net135),
    .A2(_00390_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11178_ (.A1(_04019_),
    .A2(_04020_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11179_ (.A1(_04018_),
    .A2(_04021_),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11180_ (.A1(_03957_),
    .A2(_03958_),
    .Z(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11181_ (.A1(_03957_),
    .A2(_03958_),
    .Z(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11182_ (.A1(_03956_),
    .A2(_04023_),
    .B(_04024_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11183_ (.A1(_00387_),
    .A2(_02586_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11184_ (.A1(_02762_),
    .A2(_00384_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11185_ (.A1(_02854_),
    .A2(_00381_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11186_ (.A1(_04026_),
    .A2(_04027_),
    .A3(_04028_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11187_ (.A1(_04025_),
    .A2(_04029_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11188_ (.A1(_04022_),
    .A2(_04030_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11189_ (.A1(_04015_),
    .A2(_04017_),
    .A3(_04031_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11190_ (.A1(_04012_),
    .A2(_04032_),
    .Z(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11191_ (.A1(_03981_),
    .A2(_04033_),
    .Z(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11192_ (.A1(_03979_),
    .A2(_04034_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _11193_ (.A1(_03850_),
    .A2(_03971_),
    .A3(_04035_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11194_ (.A1(_03808_),
    .A2(_03809_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11195_ (.A1(_00397_),
    .A2(_02153_),
    .A3(_03810_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11196_ (.A1(_00387_),
    .A2(_02236_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11197_ (.A1(_00381_),
    .A2(_02409_),
    .B1(_02238_),
    .B2(_00384_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11198_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02409_),
    .A4(_02238_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11199_ (.A1(_04039_),
    .A2(_04040_),
    .B(_04041_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11200_ (.I(_04042_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11201_ (.A1(_03795_),
    .A2(_03798_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11202_ (.A1(_04043_),
    .A2(_04044_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11203_ (.A1(_00397_),
    .A2(_02051_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11204_ (.A1(_00390_),
    .A2(_02236_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11205_ (.A1(_00393_),
    .A2(_02153_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11206_ (.A1(_04046_),
    .A2(_04047_),
    .A3(_04048_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11207_ (.A1(_04045_),
    .A2(_04049_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11208_ (.A1(_04043_),
    .A2(_04044_),
    .B(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11209_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02586_),
    .A4(_02584_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11210_ (.A1(_00378_),
    .A2(_02499_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11211_ (.A1(_00372_),
    .A2(_02586_),
    .B1(_02584_),
    .B2(_00375_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11212_ (.A1(_04052_),
    .A2(_04054_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11213_ (.A1(_04053_),
    .A2(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11214_ (.A1(_04052_),
    .A2(_04056_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11215_ (.A1(_00369_),
    .A2(_02762_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11216_ (.A1(_00361_),
    .A2(_02938_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11217_ (.A1(_00365_),
    .A2(_02854_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11218_ (.A1(_04059_),
    .A2(_04060_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11219_ (.A1(_04059_),
    .A2(_04060_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11220_ (.A1(_04058_),
    .A2(_04061_),
    .B(_04062_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11221_ (.A1(_03817_),
    .A2(_03820_),
    .Z(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11222_ (.A1(_04063_),
    .A2(_04064_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11223_ (.A1(_04063_),
    .A2(_04064_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11224_ (.A1(_04057_),
    .A2(_04065_),
    .B(_04066_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11225_ (.A1(_03806_),
    .A2(_03811_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11226_ (.A1(_04067_),
    .A2(_04068_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11227_ (.A1(_04067_),
    .A2(_04068_),
    .Z(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11228_ (.A1(_04051_),
    .A2(_04069_),
    .B(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11229_ (.A1(_04037_),
    .A2(_04038_),
    .B(_04071_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11230_ (.A1(_04037_),
    .A2(_04038_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11231_ (.A1(_04071_),
    .A2(_04073_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11232_ (.A1(_04051_),
    .A2(_04069_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11233_ (.A1(_04057_),
    .A2(_04065_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11234_ (.A1(_04058_),
    .A2(_04059_),
    .A3(_04060_),
    .Z(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11235_ (.A1(_00359_),
    .A2(_02938_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11236_ (.A1(net87),
    .A2(_03018_),
    .B1(_02940_),
    .B2(net84),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11237_ (.A1(net87),
    .A2(net83),
    .A3(_03018_),
    .A4(_02940_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11238_ (.A1(_04078_),
    .A2(_04079_),
    .B(_04080_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11239_ (.A1(_00351_),
    .A2(_03189_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11240_ (.A1(_00354_),
    .A2(_03018_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11241_ (.A1(_04082_),
    .A2(_04083_),
    .A3(_03855_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11242_ (.A1(_04081_),
    .A2(_04084_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11243_ (.A1(_04081_),
    .A2(_04084_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11244_ (.A1(_04077_),
    .A2(_04085_),
    .B(_04086_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11245_ (.A1(_03863_),
    .A2(_03864_),
    .Z(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11246_ (.A1(_04087_),
    .A2(_04088_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11247_ (.A1(_04087_),
    .A2(_04088_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11248_ (.A1(_04076_),
    .A2(_04089_),
    .B(_04090_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11249_ (.A1(_03866_),
    .A2(_03879_),
    .A3(_03854_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11250_ (.A1(_04091_),
    .A2(_04092_),
    .Z(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11251_ (.A1(_04076_),
    .A2(_04089_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11252_ (.A1(_04090_),
    .A2(_04094_),
    .B(_04092_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11253_ (.A1(_04075_),
    .A2(_04093_),
    .B(_04095_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11254_ (.A1(_03853_),
    .A2(_03913_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11255_ (.A1(_04096_),
    .A2(_04097_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11256_ (.A1(_04096_),
    .A2(_04097_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11257_ (.A1(_04074_),
    .A2(_04098_),
    .B(_04099_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11258_ (.A1(_03852_),
    .A2(_03969_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11259_ (.A1(_04100_),
    .A2(_04101_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11260_ (.A1(_04100_),
    .A2(_04101_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11261_ (.A1(_04072_),
    .A2(_04102_),
    .B(_04103_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11262_ (.A1(_04036_),
    .A2(_04104_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11263_ (.A1(_04072_),
    .A2(_04102_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11264_ (.A1(_00387_),
    .A2(_02153_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11265_ (.A1(_00381_),
    .A2(_02238_),
    .B1(_02236_),
    .B2(_00384_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11266_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02238_),
    .A4(_02236_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11267_ (.A1(_04107_),
    .A2(_04108_),
    .B(_04109_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11268_ (.I(_04110_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11269_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02409_),
    .A4(_02238_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11270_ (.A1(_04112_),
    .A2(_04040_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11271_ (.A1(_04039_),
    .A2(_04113_),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11272_ (.A1(_04111_),
    .A2(_04114_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11273_ (.A1(_00397_),
    .A2(_01956_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11274_ (.A1(_00390_),
    .A2(_02153_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11275_ (.A1(_00393_),
    .A2(_02051_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11276_ (.A1(_04116_),
    .A2(_04117_),
    .A3(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11277_ (.A1(_04115_),
    .A2(_04119_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11278_ (.A1(_04111_),
    .A2(_04114_),
    .B(_04120_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11279_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02584_),
    .A4(_02499_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11280_ (.A1(_00378_),
    .A2(_02409_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11281_ (.A1(_00372_),
    .A2(_02584_),
    .B1(_02499_),
    .B2(_00375_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11282_ (.A1(_04122_),
    .A2(_04124_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11283_ (.A1(_04123_),
    .A2(_04125_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11284_ (.A1(_04122_),
    .A2(_04126_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11285_ (.A1(_00369_),
    .A2(_02586_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11286_ (.A1(_00361_),
    .A2(_02854_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11287_ (.A1(_00365_),
    .A2(_02762_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11288_ (.A1(_04129_),
    .A2(_04130_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11289_ (.A1(_04129_),
    .A2(_04130_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11290_ (.A1(_04128_),
    .A2(_04131_),
    .B(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11291_ (.A1(_04053_),
    .A2(_04055_),
    .Z(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11292_ (.A1(_04133_),
    .A2(_04134_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11293_ (.A1(_04133_),
    .A2(_04134_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11294_ (.A1(_04127_),
    .A2(_04135_),
    .B(_04136_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11295_ (.A1(_04045_),
    .A2(_04049_),
    .Z(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11296_ (.A1(_04137_),
    .A2(_04138_),
    .Z(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11297_ (.A1(_04137_),
    .A2(_04138_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11298_ (.A1(_04121_),
    .A2(_04139_),
    .B(_04140_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11299_ (.A1(_04047_),
    .A2(_04048_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11300_ (.A1(_04047_),
    .A2(_04048_),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11301_ (.A1(_04046_),
    .A2(_04142_),
    .B(_04143_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11302_ (.I(_04144_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11303_ (.A1(_04141_),
    .A2(_04145_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11304_ (.A1(_04127_),
    .A2(_04135_),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11305_ (.A1(_04128_),
    .A2(_04129_),
    .A3(_04130_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11306_ (.A1(_00359_),
    .A2(_02854_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11307_ (.A1(net86),
    .A2(_02940_),
    .B1(_02938_),
    .B2(net83),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11308_ (.A1(net86),
    .A2(net83),
    .A3(_02940_),
    .A4(_02938_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11309_ (.A1(_04149_),
    .A2(_04150_),
    .B(_04151_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11310_ (.A1(_00351_),
    .A2(_03018_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11311_ (.A1(_00354_),
    .A2(_02940_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11312_ (.A1(_04153_),
    .A2(_04154_),
    .A3(_04078_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11313_ (.A1(_04152_),
    .A2(_04155_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11314_ (.A1(_04152_),
    .A2(net81),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11315_ (.A1(_04148_),
    .A2(_04156_),
    .B(_04157_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11316_ (.A1(_04077_),
    .A2(_04085_),
    .Z(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11317_ (.A1(_04158_),
    .A2(_04159_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11318_ (.A1(_04158_),
    .A2(_04159_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11319_ (.A1(_04147_),
    .A2(_04160_),
    .B(_04161_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11320_ (.A1(_04076_),
    .A2(_04089_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11321_ (.A1(_04121_),
    .A2(_04139_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11322_ (.A1(_04076_),
    .A2(_04089_),
    .A3(_04162_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _11323_ (.A1(_04094_),
    .A2(_04162_),
    .A3(_04163_),
    .B1(_04164_),
    .B2(_04165_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11324_ (.A1(_04075_),
    .A2(_04093_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11325_ (.A1(_04166_),
    .A2(_04167_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11326_ (.A1(_04166_),
    .A2(_04167_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11327_ (.A1(_04146_),
    .A2(_04168_),
    .B(_04169_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11328_ (.A1(_04074_),
    .A2(_04098_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11329_ (.A1(_04170_),
    .A2(_04171_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _11330_ (.A1(_04141_),
    .A2(_04145_),
    .A3(_04172_),
    .B1(_04171_),
    .B2(_04170_),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11331_ (.A1(_04106_),
    .A2(_04173_),
    .Z(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11332_ (.A1(_00390_),
    .A2(_00393_),
    .A3(_01249_),
    .A4(_01247_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11333_ (.A1(_00387_),
    .A2(_01247_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11334_ (.A1(_00381_),
    .A2(_01430_),
    .B1(_01249_),
    .B2(_00384_),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11335_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_01430_),
    .A4(_01249_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11336_ (.A1(_04176_),
    .A2(_04177_),
    .B(_04178_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11337_ (.I(_04179_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11338_ (.A1(_00384_),
    .A2(_01430_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11339_ (.A1(_00381_),
    .A2(_01524_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11340_ (.A1(_00387_),
    .A2(_01249_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11341_ (.A1(_04181_),
    .A2(_04182_),
    .A3(_04183_),
    .Z(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11342_ (.A1(_04180_),
    .A2(_04184_),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11343_ (.A1(_00390_),
    .A2(_01247_),
    .A3(_04185_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11344_ (.A1(_04180_),
    .A2(_04184_),
    .B(_04186_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11345_ (.A1(_00378_),
    .A2(_01524_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11346_ (.I(_04188_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11347_ (.A1(_00375_),
    .A2(_01610_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11348_ (.A1(_00372_),
    .A2(_01693_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11349_ (.A1(_04190_),
    .A2(_04191_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11350_ (.A1(_04190_),
    .A2(_04191_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11351_ (.A1(_04189_),
    .A2(_04192_),
    .B(_04193_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11352_ (.A1(_00369_),
    .A2(_01792_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11353_ (.A1(_00365_),
    .A2(_01794_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11354_ (.A1(_00361_),
    .A2(_01956_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11355_ (.A1(_04196_),
    .A2(_04197_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11356_ (.A1(_04196_),
    .A2(_04197_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11357_ (.A1(_04195_),
    .A2(_04198_),
    .B(_04199_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11358_ (.A1(_00375_),
    .A2(_01693_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11359_ (.A1(_00372_),
    .A2(_01792_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11360_ (.A1(_00378_),
    .A2(_01610_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11361_ (.I(_04203_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11362_ (.A1(_04201_),
    .A2(_04202_),
    .A3(_04204_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11363_ (.A1(_04200_),
    .A2(_04205_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11364_ (.A1(_04200_),
    .A2(_04205_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11365_ (.A1(_04194_),
    .A2(_04206_),
    .B(_04207_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11366_ (.A1(_00390_),
    .A2(_01249_),
    .B1(_01247_),
    .B2(_00393_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11367_ (.I(_04209_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11368_ (.A1(_04175_),
    .A2(_04210_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11369_ (.A1(_04181_),
    .A2(_04182_),
    .Z(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11370_ (.A1(_04181_),
    .A2(_04182_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11371_ (.A1(_04183_),
    .A2(_04212_),
    .B(_04213_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11372_ (.A1(_00384_),
    .A2(_01524_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11373_ (.A1(_00381_),
    .A2(_01610_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11374_ (.A1(_00387_),
    .A2(_01430_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11375_ (.A1(_04215_),
    .A2(_04216_),
    .A3(_04217_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11376_ (.A1(_04214_),
    .A2(_04218_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11377_ (.A1(_04211_),
    .A2(_04219_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11378_ (.A1(_04208_),
    .A2(_04220_),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11379_ (.A1(_04208_),
    .A2(_04220_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11380_ (.A1(_04187_),
    .A2(_04221_),
    .B(_04222_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11381_ (.A1(_04175_),
    .A2(_04223_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11382_ (.A1(_04175_),
    .A2(_04223_),
    .Z(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11383_ (.A1(net70),
    .A2(_01956_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11384_ (.A1(net66),
    .A2(_02153_),
    .B1(_02051_),
    .B2(net54),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11385_ (.A1(net66),
    .A2(net54),
    .A3(_02153_),
    .A4(_02051_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11386_ (.A1(_04226_),
    .A2(_04227_),
    .B(_04228_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11387_ (.A1(net83),
    .A2(_02153_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11388_ (.A1(net87),
    .A2(_02236_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11389_ (.A1(net70),
    .A2(_02051_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11390_ (.A1(_04230_),
    .A2(_04231_),
    .A3(_04232_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11391_ (.A1(_04229_),
    .A2(_04233_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11392_ (.A1(_04195_),
    .A2(_04196_),
    .A3(_04197_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11393_ (.A1(_04229_),
    .A2(_04233_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11394_ (.A1(_04234_),
    .A2(_04235_),
    .B(_04236_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11395_ (.A1(net66),
    .A2(_02236_),
    .B1(_02153_),
    .B2(net54),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11396_ (.A1(net66),
    .A2(net54),
    .A3(_02236_),
    .A4(_02153_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11397_ (.A1(_04232_),
    .A2(_04238_),
    .B(_04239_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11398_ (.A1(net84),
    .A2(_02236_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11399_ (.A1(net87),
    .A2(_02238_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11400_ (.A1(_00359_),
    .A2(_02153_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11401_ (.A1(_04241_),
    .A2(_04242_),
    .A3(_04243_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11402_ (.A1(_04240_),
    .A2(_04244_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11403_ (.A1(_00369_),
    .A2(_01794_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11404_ (.A1(_00365_),
    .A2(_01956_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11405_ (.A1(_00361_),
    .A2(_02051_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11406_ (.A1(_04246_),
    .A2(_04247_),
    .A3(_04248_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11407_ (.A1(_04245_),
    .A2(_04249_),
    .Z(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11408_ (.A1(_04237_),
    .A2(_04250_),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11409_ (.A1(_04194_),
    .A2(_04206_),
    .Z(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11410_ (.A1(_04237_),
    .A2(_04250_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11411_ (.A1(_04251_),
    .A2(_04252_),
    .B(_04253_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11412_ (.A1(_04240_),
    .A2(_04244_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11413_ (.A1(_04245_),
    .A2(_04249_),
    .B(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11414_ (.A1(net66),
    .A2(_02238_),
    .B1(_02236_),
    .B2(net54),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11415_ (.A1(net66),
    .A2(net54),
    .A3(_02238_),
    .A4(_02236_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11416_ (.A1(_04243_),
    .A2(_04257_),
    .B(_04258_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11417_ (.A1(net84),
    .A2(_02238_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11418_ (.A1(net87),
    .A2(_02409_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11419_ (.A1(_00359_),
    .A2(_02236_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11420_ (.A1(_04260_),
    .A2(_04261_),
    .A3(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11421_ (.A1(_04259_),
    .A2(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11422_ (.A1(_00369_),
    .A2(_01956_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11423_ (.A1(_00365_),
    .A2(_02051_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11424_ (.A1(_00361_),
    .A2(_02153_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11425_ (.A1(_04265_),
    .A2(_04266_),
    .A3(_04267_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11426_ (.A1(_04264_),
    .A2(_04268_),
    .Z(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11427_ (.A1(_04256_),
    .A2(_04269_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11428_ (.A1(_04201_),
    .A2(_04202_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11429_ (.A1(_04201_),
    .A2(_04202_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11430_ (.A1(_04204_),
    .A2(_04271_),
    .B(_04272_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11431_ (.A1(_04247_),
    .A2(_04248_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11432_ (.A1(_04247_),
    .A2(_04248_),
    .Z(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11433_ (.A1(_04246_),
    .A2(_04274_),
    .B(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11434_ (.A1(_00375_),
    .A2(_01792_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11435_ (.A1(_00372_),
    .A2(_01794_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11436_ (.A1(_00378_),
    .A2(_01693_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11437_ (.I(_04279_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11438_ (.A1(_04277_),
    .A2(_04278_),
    .A3(_04280_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11439_ (.A1(_04276_),
    .A2(_04281_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11440_ (.A1(_04273_),
    .A2(_04282_),
    .Z(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11441_ (.A1(_04270_),
    .A2(_04283_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11442_ (.A1(_04254_),
    .A2(_04284_),
    .Z(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11443_ (.A1(_04187_),
    .A2(_04221_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11444_ (.A1(_04251_),
    .A2(_04252_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11445_ (.A1(_04253_),
    .A2(_04287_),
    .B(_04284_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11446_ (.A1(_04285_),
    .A2(_04286_),
    .B(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11447_ (.A1(_04256_),
    .A2(_04269_),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11448_ (.A1(_04270_),
    .A2(_04283_),
    .B(_04290_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11449_ (.A1(_04259_),
    .A2(_04263_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11450_ (.A1(_04264_),
    .A2(_04268_),
    .B(_04292_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11451_ (.A1(net86),
    .A2(_02409_),
    .B1(_02238_),
    .B2(net83),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11452_ (.A1(net86),
    .A2(net83),
    .A3(_02409_),
    .A4(_02238_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11453_ (.A1(_04262_),
    .A2(_04294_),
    .B(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11454_ (.A1(_00354_),
    .A2(_02409_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11455_ (.A1(_00351_),
    .A2(_02499_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11456_ (.A1(_00359_),
    .A2(_02238_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11457_ (.A1(_04297_),
    .A2(_04298_),
    .A3(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11458_ (.A1(_04296_),
    .A2(_04300_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11459_ (.A1(_00369_),
    .A2(_02051_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11460_ (.A1(_00365_),
    .A2(_02153_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11461_ (.A1(_00361_),
    .A2(_02236_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11462_ (.A1(_04302_),
    .A2(_04303_),
    .A3(_04304_),
    .Z(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11463_ (.A1(_04301_),
    .A2(_04305_),
    .Z(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11464_ (.A1(_04293_),
    .A2(_04306_),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11465_ (.A1(_04277_),
    .A2(_04278_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11466_ (.A1(_04277_),
    .A2(_04278_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11467_ (.A1(_04280_),
    .A2(_04308_),
    .B(_04309_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11468_ (.A1(_00361_),
    .A2(_02153_),
    .B1(_02051_),
    .B2(_00365_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11469_ (.A1(_00361_),
    .A2(_00365_),
    .A3(_02153_),
    .A4(_02051_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11470_ (.A1(_04265_),
    .A2(_04311_),
    .B(_04312_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11471_ (.A1(_00375_),
    .A2(_01794_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11472_ (.A1(_00372_),
    .A2(_01956_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11473_ (.A1(_00378_),
    .A2(_01792_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11474_ (.A1(_04314_),
    .A2(_04315_),
    .A3(_04316_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11475_ (.A1(_04313_),
    .A2(_04317_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11476_ (.A1(_04310_),
    .A2(_04318_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11477_ (.A1(_04307_),
    .A2(_04319_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11478_ (.A1(_04291_),
    .A2(_04320_),
    .Z(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11479_ (.I(_04218_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11480_ (.A1(_04214_),
    .A2(_04322_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11481_ (.A1(_04211_),
    .A2(_04219_),
    .B(_04323_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11482_ (.A1(_04276_),
    .A2(_04281_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11483_ (.A1(_04273_),
    .A2(_04282_),
    .B(_04325_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11484_ (.A1(_04215_),
    .A2(_04216_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11485_ (.A1(_04215_),
    .A2(_04216_),
    .Z(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11486_ (.A1(_04217_),
    .A2(_04327_),
    .B(_04328_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11487_ (.A1(_00384_),
    .A2(_01610_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11488_ (.A1(_00381_),
    .A2(_01693_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11489_ (.A1(_00387_),
    .A2(_01524_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11490_ (.A1(_04330_),
    .A2(_04331_),
    .A3(_04332_),
    .Z(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11491_ (.A1(_04329_),
    .A2(_04333_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11492_ (.A1(_00397_),
    .A2(_01247_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11493_ (.A1(_00393_),
    .A2(_01249_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11494_ (.A1(_00390_),
    .A2(_01430_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11495_ (.A1(_04336_),
    .A2(_04337_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11496_ (.A1(_04335_),
    .A2(_04338_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11497_ (.A1(_04334_),
    .A2(_04339_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11498_ (.A1(_04324_),
    .A2(_04326_),
    .A3(_04340_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11499_ (.A1(_04321_),
    .A2(_04341_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11500_ (.A1(_04289_),
    .A2(_04342_),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11501_ (.A1(_04289_),
    .A2(_04342_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11502_ (.A1(_04225_),
    .A2(_04343_),
    .B(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11503_ (.A1(_04326_),
    .A2(_04340_),
    .Z(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11504_ (.A1(_04326_),
    .A2(_04340_),
    .Z(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11505_ (.A1(_04324_),
    .A2(_04346_),
    .B(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11506_ (.A1(_00397_),
    .A2(_01247_),
    .A3(_04338_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11507_ (.A1(_04336_),
    .A2(_04337_),
    .B(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11508_ (.I(_04350_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11509_ (.A1(_04348_),
    .A2(_04351_),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11510_ (.A1(_04270_),
    .A2(_04283_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11511_ (.A1(_04290_),
    .A2(_04353_),
    .B(_04320_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11512_ (.A1(_04321_),
    .A2(_04341_),
    .B(_04354_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11513_ (.A1(_04296_),
    .A2(_04300_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11514_ (.A1(_04301_),
    .A2(_04305_),
    .B(_04356_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11515_ (.A1(net86),
    .A2(_02499_),
    .B1(_02409_),
    .B2(net83),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11516_ (.A1(net86),
    .A2(net83),
    .A3(_02499_),
    .A4(_02409_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11517_ (.A1(_04299_),
    .A2(_04358_),
    .B(_04359_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11518_ (.A1(_00354_),
    .A2(_02499_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11519_ (.A1(_00351_),
    .A2(_02584_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11520_ (.A1(_00359_),
    .A2(_02409_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11521_ (.A1(_04361_),
    .A2(_04362_),
    .A3(_04363_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11522_ (.A1(_04364_),
    .A2(_04360_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11523_ (.A1(_00369_),
    .A2(_02153_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11524_ (.A1(_00365_),
    .A2(_02236_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11525_ (.A1(_00361_),
    .A2(_02238_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11526_ (.A1(_04366_),
    .A2(_04367_),
    .A3(_04368_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11527_ (.A1(_04369_),
    .A2(_04365_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11528_ (.A1(_04357_),
    .A2(_04370_),
    .Z(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11529_ (.I(_04316_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11530_ (.A1(_04314_),
    .A2(_04315_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11531_ (.A1(_04314_),
    .A2(_04315_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11532_ (.A1(_04372_),
    .A2(_04373_),
    .B(_04374_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11533_ (.A1(_04303_),
    .A2(_04304_),
    .Z(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11534_ (.A1(_04303_),
    .A2(_04304_),
    .Z(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11535_ (.A1(_04302_),
    .A2(_04376_),
    .B(_04377_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11536_ (.A1(_00375_),
    .A2(_01956_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11537_ (.A1(_00372_),
    .A2(_02051_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11538_ (.A1(_00378_),
    .A2(_01794_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11539_ (.I(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11540_ (.A1(_04379_),
    .A2(_04380_),
    .A3(_04382_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11541_ (.A1(_04378_),
    .A2(_04383_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11542_ (.A1(_04375_),
    .A2(_04384_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11543_ (.A1(_04293_),
    .A2(_04306_),
    .Z(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11544_ (.A1(_04307_),
    .A2(_04319_),
    .B(_04386_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11545_ (.A1(_04371_),
    .A2(_04385_),
    .A3(_04387_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11546_ (.I(_04333_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11547_ (.A1(_04329_),
    .A2(_04389_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11548_ (.A1(_04334_),
    .A2(_04339_),
    .B(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11549_ (.A1(_04313_),
    .A2(_04317_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11550_ (.A1(_04310_),
    .A2(_04318_),
    .B(_04392_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11551_ (.A1(_00381_),
    .A2(_01693_),
    .B1(_01610_),
    .B2(_00384_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11552_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_01693_),
    .A4(_01610_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11553_ (.A1(_04332_),
    .A2(_04394_),
    .B(_04395_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11554_ (.A1(_00384_),
    .A2(_01693_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11555_ (.A1(_00381_),
    .A2(_01792_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11556_ (.A1(_00387_),
    .A2(_01610_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11557_ (.A1(_04397_),
    .A2(_04398_),
    .A3(_04399_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11558_ (.A1(_04396_),
    .A2(_04400_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11559_ (.A1(_00397_),
    .A2(_01249_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11560_ (.A1(_00393_),
    .A2(_01430_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11561_ (.A1(_00390_),
    .A2(_01524_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11562_ (.A1(_04403_),
    .A2(_04404_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11563_ (.A1(_04402_),
    .A2(_04405_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11564_ (.A1(_04401_),
    .A2(_04406_),
    .Z(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11565_ (.A1(_04391_),
    .A2(_04393_),
    .A3(_04407_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11566_ (.A1(_04388_),
    .A2(_04408_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11567_ (.A1(_04409_),
    .A2(_04355_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11568_ (.A1(_04352_),
    .A2(_04410_),
    .Z(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11569_ (.A1(_04345_),
    .A2(_04411_),
    .Z(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11570_ (.A1(_04224_),
    .A2(_04412_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11571_ (.A1(_00381_),
    .A2(_01249_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11572_ (.A1(_00384_),
    .A2(_01247_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11573_ (.A1(_04414_),
    .A2(_04415_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11574_ (.A1(_00381_),
    .A2(_01430_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11575_ (.A1(_00384_),
    .A2(_01249_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11576_ (.A1(_04417_),
    .A2(_04418_),
    .A3(_04176_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11577_ (.A1(_04416_),
    .A2(_04419_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11578_ (.A1(_00378_),
    .A2(_01430_),
    .Z(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11579_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_01610_),
    .A4(_01524_),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11580_ (.A1(_00372_),
    .A2(_01610_),
    .B1(_01524_),
    .B2(_00375_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11581_ (.A1(_04422_),
    .A2(_04423_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11582_ (.A1(_04421_),
    .A2(_04424_),
    .B(_04422_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11583_ (.A1(_00369_),
    .A2(_01693_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11584_ (.A1(_00365_),
    .A2(_01792_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11585_ (.A1(_00361_),
    .A2(_01794_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11586_ (.A1(_04427_),
    .A2(_04428_),
    .Z(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11587_ (.A1(_04427_),
    .A2(_04428_),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11588_ (.A1(_04426_),
    .A2(_04429_),
    .B(_04430_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11589_ (.A1(_04190_),
    .A2(_04191_),
    .A3(_04189_),
    .Z(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11590_ (.A1(_04431_),
    .A2(_04432_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11591_ (.A1(_04431_),
    .A2(_04432_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11592_ (.A1(_04425_),
    .A2(_04433_),
    .B(_04434_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11593_ (.A1(_00390_),
    .A2(_01247_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11594_ (.A1(_04436_),
    .A2(_04185_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11595_ (.A1(_04435_),
    .A2(_04437_),
    .Z(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11596_ (.A1(_04435_),
    .A2(_04437_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11597_ (.A1(_04420_),
    .A2(_04438_),
    .B(_04439_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11598_ (.A1(_04425_),
    .A2(_04433_),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11599_ (.A1(_04426_),
    .A2(_04427_),
    .A3(_04428_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11600_ (.A1(net70),
    .A2(_01794_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11601_ (.A1(net66),
    .A2(_02051_),
    .B1(_01956_),
    .B2(net54),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11602_ (.A1(net66),
    .A2(net54),
    .A3(_02051_),
    .A4(_01956_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11603_ (.A1(_04443_),
    .A2(_04444_),
    .B(_04445_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11604_ (.A1(net54),
    .A2(_02051_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11605_ (.A1(net86),
    .A2(_02153_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11606_ (.A1(_04447_),
    .A2(_04448_),
    .A3(_04226_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11607_ (.A1(_04446_),
    .A2(_04449_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11608_ (.A1(_04446_),
    .A2(_04449_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11609_ (.A1(_04442_),
    .A2(_04450_),
    .B(_04451_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11610_ (.A1(_04234_),
    .A2(_04235_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11611_ (.A1(_04452_),
    .A2(_04453_),
    .Z(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11612_ (.A1(_04452_),
    .A2(_04453_),
    .Z(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11613_ (.A1(_04441_),
    .A2(_04454_),
    .B(_04455_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11614_ (.A1(_04251_),
    .A2(_04252_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11615_ (.A1(_04420_),
    .A2(_04435_),
    .A3(_04437_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11616_ (.A1(_04251_),
    .A2(_04252_),
    .A3(_04456_),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _11617_ (.A1(_04287_),
    .A2(_04456_),
    .A3(_04457_),
    .B1(_04458_),
    .B2(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11618_ (.A1(_04285_),
    .A2(_04286_),
    .Z(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11619_ (.A1(_04460_),
    .A2(_04461_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11620_ (.A1(_04460_),
    .A2(_04461_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _11621_ (.A1(_04440_),
    .A2(_04462_),
    .B(_04463_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _11622_ (.A1(_04289_),
    .A2(_04342_),
    .A3(_04225_),
    .Z(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11623_ (.A1(_04464_),
    .A2(_04465_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11624_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_01524_),
    .A4(_01430_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11625_ (.A1(_00378_),
    .A2(_01249_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11626_ (.A1(_00372_),
    .A2(_01524_),
    .B1(_01430_),
    .B2(_00375_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11627_ (.A1(_04467_),
    .A2(_04469_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11628_ (.A1(_04468_),
    .A2(_04470_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11629_ (.A1(_04467_),
    .A2(_04471_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11630_ (.A1(_00361_),
    .A2(_00365_),
    .A3(_01792_),
    .A4(_01693_),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11631_ (.A1(_00369_),
    .A2(_01610_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11632_ (.A1(_00361_),
    .A2(_01792_),
    .B1(_01693_),
    .B2(_00365_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11633_ (.A1(_04474_),
    .A2(_04473_),
    .A3(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11634_ (.A1(_04473_),
    .A2(_04476_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11635_ (.A1(_04421_),
    .A2(_04424_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11636_ (.A1(_04477_),
    .A2(_04478_),
    .Z(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11637_ (.I(_04478_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11638_ (.A1(_04477_),
    .A2(_04480_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11639_ (.A1(_04472_),
    .A2(_04479_),
    .B(_04481_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11640_ (.A1(_04416_),
    .A2(_04419_),
    .Z(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11641_ (.A1(_04482_),
    .A2(_04483_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11642_ (.A1(net70),
    .A2(_01792_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11643_ (.A1(net66),
    .A2(_01956_),
    .B1(_01794_),
    .B2(net54),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11644_ (.A1(net66),
    .A2(net54),
    .A3(_01956_),
    .A4(_01794_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11645_ (.A1(_04485_),
    .A2(_04486_),
    .B(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11646_ (.A1(net54),
    .A2(_01956_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11647_ (.A1(net66),
    .A2(_02051_),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11648_ (.A1(_04489_),
    .A2(_04490_),
    .A3(_04443_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11649_ (.A1(_04488_),
    .A2(_04491_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11650_ (.A1(_04473_),
    .A2(_04475_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11651_ (.A1(_04474_),
    .A2(_04493_),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11652_ (.A1(_04488_),
    .A2(_04491_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11653_ (.A1(_04492_),
    .A2(_04494_),
    .B(_04495_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11654_ (.A1(_04442_),
    .A2(_04450_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11655_ (.A1(_04496_),
    .A2(_04497_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11656_ (.A1(_04472_),
    .A2(_04479_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11657_ (.A1(_04496_),
    .A2(_04497_),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11658_ (.A1(_04498_),
    .A2(_04499_),
    .B(_04500_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11659_ (.A1(_04441_),
    .A2(_04454_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11660_ (.A1(_04501_),
    .A2(_04502_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11661_ (.A1(_04501_),
    .A2(_04502_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11662_ (.A1(_04484_),
    .A2(_04503_),
    .B(_04504_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11663_ (.A1(_04458_),
    .A2(_04459_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11664_ (.A1(_04505_),
    .A2(_04506_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11665_ (.A1(_04482_),
    .A2(_04483_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11666_ (.I(_04508_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11667_ (.A1(_04505_),
    .A2(_04506_),
    .Z(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11668_ (.A1(_04509_),
    .A2(_04510_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11669_ (.A1(_04460_),
    .A2(_04461_),
    .A3(_04440_),
    .Z(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11670_ (.A1(_04507_),
    .A2(_04511_),
    .B(_04512_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11671_ (.A1(_04464_),
    .A2(_04465_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11672_ (.A1(_04513_),
    .A2(_04514_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11673_ (.A1(_04466_),
    .A2(_04515_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11674_ (.A1(_04505_),
    .A2(_04506_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11675_ (.A1(_04508_),
    .A2(_04517_),
    .B(_04507_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11676_ (.A1(_04518_),
    .A2(_04512_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11677_ (.I(_04519_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11678_ (.A1(_00361_),
    .A2(_00365_),
    .A3(_01610_),
    .A4(_01524_),
    .Z(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11679_ (.A1(_00369_),
    .A2(_01430_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11680_ (.A1(_00361_),
    .A2(_01610_),
    .B1(_01524_),
    .B2(_00365_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11681_ (.A1(_04522_),
    .A2(_04521_),
    .A3(_04523_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11682_ (.A1(_04521_),
    .A2(_04524_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11683_ (.A1(_00378_),
    .A2(_01247_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11684_ (.A1(_00372_),
    .A2(_01430_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11685_ (.A1(_00375_),
    .A2(_01249_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11686_ (.A1(_04527_),
    .A2(_04528_),
    .Z(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11687_ (.A1(_04526_),
    .A2(_04529_),
    .Z(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11688_ (.A1(_00372_),
    .A2(_01249_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11689_ (.A1(_00375_),
    .A2(_01247_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11690_ (.A1(_04531_),
    .A2(_04532_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11691_ (.I(_04533_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11692_ (.A1(_04525_),
    .A2(_04530_),
    .Z(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11693_ (.A1(_04534_),
    .A2(_04535_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11694_ (.A1(_04525_),
    .A2(_04530_),
    .B(_04536_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11695_ (.A1(_00381_),
    .A2(_01247_),
    .A3(_04537_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11696_ (.A1(_00381_),
    .A2(_01247_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11697_ (.A1(_04539_),
    .A2(_04537_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11698_ (.A1(net70),
    .A2(_01610_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11699_ (.A1(net66),
    .A2(_01792_),
    .B1(_01693_),
    .B2(net54),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11700_ (.A1(net66),
    .A2(net54),
    .A3(_01792_),
    .A4(_01693_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11701_ (.A1(_04541_),
    .A2(_04542_),
    .B(_04543_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11702_ (.A1(net86),
    .A2(_01794_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11703_ (.A1(net54),
    .A2(_01792_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11704_ (.A1(net70),
    .A2(_01693_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11705_ (.A1(_04545_),
    .A2(_04546_),
    .A3(_04547_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11706_ (.A1(_04544_),
    .A2(_04548_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11707_ (.A1(_04521_),
    .A2(_04523_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11708_ (.A1(_04522_),
    .A2(_04550_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11709_ (.A1(_04544_),
    .A2(_04548_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11710_ (.A1(_04549_),
    .A2(_04551_),
    .B(_04552_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11711_ (.A1(net66),
    .A2(_01794_),
    .B1(_01792_),
    .B2(net54),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11712_ (.A1(net66),
    .A2(net54),
    .A3(_01794_),
    .A4(_01792_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11713_ (.A1(_04547_),
    .A2(_04554_),
    .B(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11714_ (.A1(net66),
    .A2(_01956_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11715_ (.A1(net54),
    .A2(_01794_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11716_ (.A1(_04557_),
    .A2(_04558_),
    .A3(_04485_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11717_ (.A1(_04556_),
    .A2(_04559_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11718_ (.A1(_00369_),
    .A2(_01524_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11719_ (.A1(_00361_),
    .A2(_00365_),
    .A3(_01693_),
    .A4(_01610_),
    .Z(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11720_ (.A1(_00361_),
    .A2(_01693_),
    .B1(_01610_),
    .B2(_00365_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11721_ (.A1(_04562_),
    .A2(_04563_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11722_ (.A1(_04561_),
    .A2(_04564_),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11723_ (.A1(_04560_),
    .A2(_04565_),
    .Z(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11724_ (.A1(_04553_),
    .A2(_04566_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11725_ (.A1(_04533_),
    .A2(_04535_),
    .Z(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11726_ (.A1(_04553_),
    .A2(_04566_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11727_ (.A1(_04567_),
    .A2(_04568_),
    .B(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11728_ (.A1(_04556_),
    .A2(_04559_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11729_ (.A1(_04560_),
    .A2(_04565_),
    .B(_04571_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11730_ (.A1(_04492_),
    .A2(_04494_),
    .Z(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11731_ (.A1(_04572_),
    .A2(_04573_),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11732_ (.A1(_00378_),
    .A2(_01247_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11733_ (.A1(_04527_),
    .A2(_04528_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11734_ (.A1(_04575_),
    .A2(_04529_),
    .B(_04576_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11735_ (.A1(_04561_),
    .A2(_04562_),
    .A3(_04563_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11736_ (.A1(_04562_),
    .A2(_04578_),
    .Z(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11737_ (.A1(_04468_),
    .A2(_04470_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11738_ (.A1(_04579_),
    .A2(_04580_),
    .Z(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11739_ (.A1(_04577_),
    .A2(_04581_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11740_ (.A1(_04574_),
    .A2(_04582_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11741_ (.A1(_04570_),
    .A2(_04583_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11742_ (.A1(_04570_),
    .A2(_04583_),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11743_ (.A1(_04540_),
    .A2(_04584_),
    .B(_04585_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11744_ (.I(_04580_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11745_ (.A1(_04579_),
    .A2(_04587_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11746_ (.A1(_04577_),
    .A2(_04581_),
    .B(_04588_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11747_ (.A1(_04414_),
    .A2(_04415_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11748_ (.A1(_04416_),
    .A2(_04590_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11749_ (.A1(_04589_),
    .A2(_04591_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11750_ (.A1(_04572_),
    .A2(_04573_),
    .Z(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11751_ (.A1(_04574_),
    .A2(_04582_),
    .B(_04593_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11752_ (.A1(_04498_),
    .A2(_04499_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11753_ (.A1(_04594_),
    .A2(_04595_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11754_ (.A1(_04592_),
    .A2(_04596_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11755_ (.A1(_04586_),
    .A2(_04597_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11756_ (.A1(_04586_),
    .A2(_04597_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11757_ (.A1(_04538_),
    .A2(_04598_),
    .B(_04599_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11758_ (.A1(_04416_),
    .A2(_04589_),
    .A3(_04590_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11759_ (.A1(_04594_),
    .A2(_04595_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11760_ (.A1(_04592_),
    .A2(_04596_),
    .B(_04602_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11761_ (.A1(_04484_),
    .A2(_04503_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11762_ (.A1(_04601_),
    .A2(_04603_),
    .A3(_04604_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11763_ (.A1(_04600_),
    .A2(_04605_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11764_ (.A1(_04603_),
    .A2(_04604_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11765_ (.A1(_04603_),
    .A2(_04604_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11766_ (.A1(_04601_),
    .A2(_04607_),
    .B(_04608_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11767_ (.A1(_04509_),
    .A2(_04510_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11768_ (.A1(_04609_),
    .A2(_04610_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11769_ (.A1(_04609_),
    .A2(_04610_),
    .Z(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11770_ (.A1(_04606_),
    .A2(_04611_),
    .B(_04612_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11771_ (.A1(_04570_),
    .A2(_04583_),
    .A3(_04540_),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11772_ (.A1(_00361_),
    .A2(_00365_),
    .A3(_01524_),
    .A4(_01430_),
    .Z(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11773_ (.A1(_00361_),
    .A2(_01524_),
    .B1(_01430_),
    .B2(_00365_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11774_ (.A1(_04615_),
    .A2(_04616_),
    .Z(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11775_ (.A1(_00369_),
    .A2(_01249_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11776_ (.A1(_04617_),
    .A2(_04618_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11777_ (.A1(_04615_),
    .A2(_04619_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11778_ (.A1(_04531_),
    .A2(_04532_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11779_ (.A1(_04533_),
    .A2(_04621_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11780_ (.A1(_04620_),
    .A2(_04622_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11781_ (.A1(_04620_),
    .A2(_04622_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11782_ (.A1(net70),
    .A2(_01524_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11783_ (.A1(net66),
    .A2(_01693_),
    .B1(_01610_),
    .B2(net54),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11784_ (.A1(net66),
    .A2(net54),
    .A3(_01693_),
    .A4(_01610_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11785_ (.A1(_04625_),
    .A2(_04626_),
    .B(_04627_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11786_ (.A1(net66),
    .A2(_01792_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11787_ (.A1(net54),
    .A2(_01693_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11788_ (.A1(_04629_),
    .A2(_04630_),
    .A3(_04541_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11789_ (.A1(_04628_),
    .A2(_04631_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11790_ (.A1(_04617_),
    .A2(_04618_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11791_ (.A1(_04628_),
    .A2(_04631_),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11792_ (.A1(_04632_),
    .A2(_04633_),
    .B(_04634_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11793_ (.A1(_04549_),
    .A2(_04551_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11794_ (.A1(_04635_),
    .A2(_04636_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11795_ (.A1(_04635_),
    .A2(_04636_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11796_ (.A1(_04624_),
    .A2(_04637_),
    .B(_04638_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11797_ (.A1(_04553_),
    .A2(_04566_),
    .A3(_04568_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11798_ (.A1(_04639_),
    .A2(_04640_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11799_ (.A1(_04639_),
    .A2(_04640_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11800_ (.A1(_04623_),
    .A2(_04641_),
    .B(_04642_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _11801_ (.A1(_04614_),
    .A2(_04643_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11802_ (.A1(_04623_),
    .A2(_04639_),
    .A3(_04640_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11803_ (.A1(_00361_),
    .A2(_00365_),
    .A3(_01430_),
    .A4(_01249_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11804_ (.A1(_00369_),
    .A2(_01247_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11805_ (.A1(_00361_),
    .A2(_01430_),
    .B1(_01249_),
    .B2(_00365_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11806_ (.A1(_04647_),
    .A2(_04646_),
    .A3(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11807_ (.A1(_04646_),
    .A2(_04649_),
    .Z(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11808_ (.A1(_00372_),
    .A2(_01247_),
    .A3(_04650_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11809_ (.A1(_00372_),
    .A2(_01247_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11810_ (.A1(_04652_),
    .A2(_04650_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11811_ (.I(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11812_ (.A1(_04646_),
    .A2(_04648_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11813_ (.A1(_04647_),
    .A2(_04655_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11814_ (.A1(net70),
    .A2(_01430_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11815_ (.A1(net66),
    .A2(_01610_),
    .B1(_01524_),
    .B2(net54),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11816_ (.A1(net66),
    .A2(net54),
    .A3(_01610_),
    .A4(_01524_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11817_ (.A1(_04657_),
    .A2(_04658_),
    .B(_04659_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11818_ (.A1(net66),
    .A2(_01693_),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11819_ (.A1(net54),
    .A2(_01610_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11820_ (.A1(_04661_),
    .A2(_04662_),
    .A3(_04625_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11821_ (.A1(_04660_),
    .A2(_04663_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11822_ (.A1(_04660_),
    .A2(_04663_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11823_ (.A1(_04656_),
    .A2(_04664_),
    .B(_04665_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11824_ (.A1(_04632_),
    .A2(_04633_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11825_ (.A1(_04666_),
    .A2(_04667_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11826_ (.A1(_04666_),
    .A2(_04667_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11827_ (.A1(_04654_),
    .A2(_04668_),
    .B(_04669_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11828_ (.A1(_04635_),
    .A2(_04636_),
    .A3(_04624_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11829_ (.A1(_04670_),
    .A2(_04671_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11830_ (.A1(_04670_),
    .A2(_04671_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11831_ (.A1(_04651_),
    .A2(_04672_),
    .B(_04673_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11832_ (.A1(_04645_),
    .A2(_04674_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11833_ (.A1(_00361_),
    .A2(_00365_),
    .A3(_01249_),
    .A4(_01247_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11834_ (.A1(_00361_),
    .A2(_01249_),
    .B1(_01247_),
    .B2(_00365_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11835_ (.I(_04677_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11836_ (.A1(_04676_),
    .A2(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11837_ (.A1(net70),
    .A2(_01249_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11838_ (.A1(net66),
    .A2(_01524_),
    .B1(_01430_),
    .B2(net54),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11839_ (.A1(net66),
    .A2(net54),
    .A3(_01524_),
    .A4(_01430_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11840_ (.A1(_04680_),
    .A2(_04681_),
    .B(_04682_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11841_ (.A1(net66),
    .A2(_01610_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11842_ (.A1(net54),
    .A2(_01524_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11843_ (.A1(net70),
    .A2(_01430_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11844_ (.A1(_04684_),
    .A2(_04685_),
    .A3(_04686_),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11845_ (.A1(_04683_),
    .A2(_04687_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11846_ (.A1(_04683_),
    .A2(_04687_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11847_ (.A1(_04679_),
    .A2(_04688_),
    .B(_04689_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11848_ (.A1(_04656_),
    .A2(_04664_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11849_ (.A1(_04690_),
    .A2(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11850_ (.A1(_04690_),
    .A2(_04691_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11851_ (.A1(_04676_),
    .A2(_04692_),
    .B(_04693_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _11852_ (.A1(_04666_),
    .A2(_04667_),
    .A3(_04653_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11853_ (.A1(_04651_),
    .A2(_04670_),
    .A3(_04671_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11854_ (.A1(_04694_),
    .A2(_04695_),
    .A3(_04696_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11855_ (.A1(_04645_),
    .A2(_04674_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11856_ (.A1(_04675_),
    .A2(_04697_),
    .B(_04698_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11857_ (.A1(_04644_),
    .A2(_04699_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11858_ (.A1(_04676_),
    .A2(_04690_),
    .A3(_04691_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11859_ (.A1(_04694_),
    .A2(_04695_),
    .B(_04701_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11860_ (.A1(_04694_),
    .A2(_04695_),
    .B(_04696_),
    .C(_04702_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11861_ (.A1(_04645_),
    .A2(_04674_),
    .A3(_04697_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11862_ (.A1(net66),
    .A2(_01524_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11863_ (.A1(net54),
    .A2(_01430_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11864_ (.A1(_04705_),
    .A2(_04706_),
    .A3(_04680_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11865_ (.A1(net66),
    .A2(_01430_),
    .B1(_01249_),
    .B2(net54),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11866_ (.A1(net70),
    .A2(_01247_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11867_ (.A1(net66),
    .A2(net54),
    .A3(_01430_),
    .A4(_01249_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11868_ (.A1(_04708_),
    .A2(_04709_),
    .B(_04710_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11869_ (.A1(_04707_),
    .A2(_04711_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11870_ (.A1(_04707_),
    .A2(_04711_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11871_ (.A1(_00361_),
    .A2(_01247_),
    .A3(_04713_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11872_ (.A1(_04712_),
    .A2(_04714_),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11873_ (.A1(_04679_),
    .A2(_04688_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11874_ (.A1(_04715_),
    .A2(_04716_),
    .Z(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11875_ (.A1(_04717_),
    .A2(_04703_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11876_ (.A1(_04704_),
    .A2(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11877_ (.A1(net70),
    .A2(_01430_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11878_ (.A1(net66),
    .A2(net54),
    .A3(_01249_),
    .A4(_01247_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11879_ (.A1(_04686_),
    .A2(_04720_),
    .B(_04721_),
    .C(_04714_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11880_ (.A1(_00361_),
    .A2(_01247_),
    .B(_04713_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11881_ (.A1(_04722_),
    .A2(_04723_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11882_ (.A1(_04715_),
    .A2(_04716_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11883_ (.A1(_04717_),
    .A2(_04724_),
    .A3(_04725_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11884_ (.A1(_04704_),
    .A2(_04718_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11885_ (.A1(_04703_),
    .A2(_04719_),
    .A3(_04726_),
    .B(_04727_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11886_ (.A1(_04614_),
    .A2(_04643_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _11887_ (.A1(_04644_),
    .A2(_04698_),
    .B(_04729_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11888_ (.A1(_04538_),
    .A2(_04598_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11889_ (.A1(_04644_),
    .A2(_04675_),
    .A3(_04697_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11890_ (.A1(_04700_),
    .A2(_04728_),
    .B1(_04730_),
    .B2(_04731_),
    .C(_04732_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11891_ (.A1(_04600_),
    .A2(_04605_),
    .Z(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11892_ (.A1(_04730_),
    .A2(_04731_),
    .B(_04734_),
    .C(_04611_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _11893_ (.A1(_04520_),
    .A2(_04613_),
    .B1(_04733_),
    .B2(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11894_ (.A1(_04519_),
    .A2(_04612_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11895_ (.A1(_04513_),
    .A2(_04514_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11896_ (.A1(_04737_),
    .A2(_04738_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _11897_ (.A1(_04413_),
    .A2(_04516_),
    .B1(_04736_),
    .B2(_04739_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11898_ (.A1(_04464_),
    .A2(_04465_),
    .B(_04413_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _11899_ (.A1(_04741_),
    .A2(_04740_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11900_ (.A1(_00387_),
    .A2(_01956_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11901_ (.A1(_00381_),
    .A2(_02153_),
    .B1(_02051_),
    .B2(_00384_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11902_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02153_),
    .A4(_02051_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11903_ (.A1(_04743_),
    .A2(_04744_),
    .B(_04745_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11904_ (.I(_04746_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11905_ (.A1(_00387_),
    .A2(_02051_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11906_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02236_),
    .A4(_02153_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11907_ (.A1(_00381_),
    .A2(_02236_),
    .B1(_02153_),
    .B2(_00384_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11908_ (.A1(_04749_),
    .A2(_04750_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11909_ (.A1(_04748_),
    .A2(_04751_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11910_ (.A1(_04747_),
    .A2(_04752_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11911_ (.A1(_00397_),
    .A2(_01792_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11912_ (.A1(_00390_),
    .A2(_01956_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11913_ (.A1(_00393_),
    .A2(_01794_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11914_ (.A1(_04754_),
    .A2(_04755_),
    .A3(_04756_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11915_ (.A1(_04753_),
    .A2(_04757_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11916_ (.A1(_04747_),
    .A2(_04752_),
    .B(_04758_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11917_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02409_),
    .A4(_02238_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11918_ (.A1(_00378_),
    .A2(_02236_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11919_ (.A1(_00372_),
    .A2(_02409_),
    .B1(_02238_),
    .B2(_00375_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11920_ (.A1(_04760_),
    .A2(_04762_),
    .Z(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11921_ (.A1(_04761_),
    .A2(_04763_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11922_ (.A1(_04760_),
    .A2(_04764_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11923_ (.A1(_00369_),
    .A2(_02499_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11924_ (.A1(_00361_),
    .A2(_02586_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11925_ (.A1(_00365_),
    .A2(net135),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11926_ (.A1(_04767_),
    .A2(_04768_),
    .Z(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11927_ (.A1(_04767_),
    .A2(_04768_),
    .Z(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11928_ (.A1(_04766_),
    .A2(_04769_),
    .B(_04770_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11929_ (.A1(_00378_),
    .A2(_02238_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11930_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02499_),
    .A4(_02409_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11931_ (.A1(_00372_),
    .A2(_02499_),
    .B1(_02409_),
    .B2(_00375_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11932_ (.A1(_04773_),
    .A2(_04774_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11933_ (.A1(_04772_),
    .A2(_04775_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11934_ (.A1(_04771_),
    .A2(_04776_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11935_ (.A1(_04771_),
    .A2(_04776_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11936_ (.A1(_04765_),
    .A2(_04777_),
    .B(_04778_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11937_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02236_),
    .A4(_02153_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11938_ (.A1(_04748_),
    .A2(_04750_),
    .B(_04780_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11939_ (.I(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11940_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02238_),
    .A4(_02236_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11941_ (.A1(_04783_),
    .A2(_04108_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11942_ (.A1(_04107_),
    .A2(_04784_),
    .Z(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11943_ (.A1(_04782_),
    .A2(_04785_),
    .Z(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11944_ (.A1(_00397_),
    .A2(_01794_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11945_ (.A1(_00390_),
    .A2(_02051_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11946_ (.A1(_00393_),
    .A2(_01956_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11947_ (.A1(_04787_),
    .A2(_04788_),
    .A3(_04789_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11948_ (.A1(_04786_),
    .A2(_04790_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11949_ (.A1(_04779_),
    .A2(_04791_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11950_ (.A1(_04779_),
    .A2(_04791_),
    .Z(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11951_ (.A1(_04759_),
    .A2(_04792_),
    .B(_04793_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11952_ (.A1(_04788_),
    .A2(_04789_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11953_ (.A1(_04788_),
    .A2(_04789_),
    .Z(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11954_ (.A1(_04787_),
    .A2(_04795_),
    .B(_04796_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11955_ (.I(_04797_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11956_ (.A1(_04794_),
    .A2(_04798_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11957_ (.I(_04799_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11958_ (.A1(_04794_),
    .A2(_04797_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11959_ (.A1(_04759_),
    .A2(_04792_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11960_ (.A1(_04765_),
    .A2(_04777_),
    .Z(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11961_ (.A1(_04766_),
    .A2(_04767_),
    .A3(_04768_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11962_ (.A1(_00359_),
    .A2(_02586_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11963_ (.A1(net66),
    .A2(_02854_),
    .B1(_02762_),
    .B2(net83),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11964_ (.A1(net66),
    .A2(net83),
    .A3(_02854_),
    .A4(_02762_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11965_ (.A1(_04805_),
    .A2(_04806_),
    .B(_04807_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11966_ (.A1(_00351_),
    .A2(_02938_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11967_ (.A1(_00354_),
    .A2(_02854_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11968_ (.A1(_00359_),
    .A2(_02762_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11969_ (.A1(_04809_),
    .A2(_04810_),
    .A3(_04811_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11970_ (.A1(_04808_),
    .A2(_04812_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11971_ (.A1(_04808_),
    .A2(_04812_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11972_ (.A1(_04804_),
    .A2(_04813_),
    .B(_04814_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11973_ (.A1(_00369_),
    .A2(_02584_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11974_ (.A1(_00361_),
    .A2(_02762_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11975_ (.A1(_00365_),
    .A2(_02586_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _11976_ (.A1(_04816_),
    .A2(_04817_),
    .A3(_04818_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11977_ (.A1(net86),
    .A2(_02938_),
    .B1(_02854_),
    .B2(net83),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11978_ (.A1(net86),
    .A2(net83),
    .A3(_02938_),
    .A4(_02854_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11979_ (.A1(_04811_),
    .A2(_04820_),
    .B(_04821_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11980_ (.A1(_00351_),
    .A2(_02940_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11981_ (.A1(_00354_),
    .A2(_02938_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11982_ (.A1(_04823_),
    .A2(_04824_),
    .A3(_04149_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11983_ (.A1(_04822_),
    .A2(_04825_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11984_ (.A1(_04819_),
    .A2(_04826_),
    .Z(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11985_ (.A1(_04815_),
    .A2(_04827_),
    .Z(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11986_ (.A1(_04815_),
    .A2(_04827_),
    .Z(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11987_ (.A1(_04803_),
    .A2(_04828_),
    .B(_04829_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11988_ (.A1(_04772_),
    .A2(_04775_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11989_ (.A1(_04773_),
    .A2(_04831_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11990_ (.A1(_04817_),
    .A2(_04818_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11991_ (.A1(_04817_),
    .A2(_04818_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11992_ (.A1(_04816_),
    .A2(_04833_),
    .B(_04834_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11993_ (.A1(_04123_),
    .A2(_04125_),
    .Z(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11994_ (.A1(_04835_),
    .A2(_04836_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11995_ (.A1(_04832_),
    .A2(_04837_),
    .Z(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11996_ (.A1(_04822_),
    .A2(_04825_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11997_ (.A1(_04819_),
    .A2(_04826_),
    .B(_04839_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11998_ (.A1(_04148_),
    .A2(_04156_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11999_ (.A1(_04840_),
    .A2(_04841_),
    .Z(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12000_ (.A1(_04838_),
    .A2(_04842_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12001_ (.A1(_04830_),
    .A2(_04843_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12002_ (.A1(_04830_),
    .A2(_04843_),
    .Z(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12003_ (.A1(_04802_),
    .A2(_04844_),
    .B(_04845_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12004_ (.A1(_04786_),
    .A2(_04790_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12005_ (.A1(_04782_),
    .A2(_04785_),
    .B(_04847_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12006_ (.A1(_04835_),
    .A2(_04836_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12007_ (.A1(_04832_),
    .A2(_04837_),
    .B(_04849_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12008_ (.A1(_04115_),
    .A2(_04119_),
    .Z(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12009_ (.A1(_04850_),
    .A2(_04851_),
    .Z(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12010_ (.A1(_04852_),
    .A2(_04848_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12011_ (.A1(_04840_),
    .A2(_04841_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12012_ (.A1(_04838_),
    .A2(_04842_),
    .B(_04854_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12013_ (.A1(_04147_),
    .A2(_04160_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12014_ (.A1(_04855_),
    .A2(_04856_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12015_ (.A1(_04853_),
    .A2(_04857_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12016_ (.A1(_04858_),
    .A2(_04846_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12017_ (.A1(_04846_),
    .A2(_04858_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12018_ (.A1(_04801_),
    .A2(net99),
    .B(_04860_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12019_ (.A1(_04855_),
    .A2(_04856_),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12020_ (.A1(net89),
    .A2(_04857_),
    .B(_04862_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12021_ (.A1(_04164_),
    .A2(_04165_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12022_ (.A1(_04850_),
    .A2(_04851_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12023_ (.A1(_04848_),
    .A2(_04852_),
    .B(_04865_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12024_ (.A1(_04117_),
    .A2(_04118_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12025_ (.A1(_04117_),
    .A2(_04118_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12026_ (.A1(_04116_),
    .A2(_04867_),
    .B(_04868_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12027_ (.A1(_04866_),
    .A2(_04869_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12028_ (.A1(_04863_),
    .A2(_04864_),
    .A3(_04870_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12029_ (.A1(_04800_),
    .A2(_04861_),
    .A3(_04871_),
    .Z(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12030_ (.A1(_00387_),
    .A2(_01794_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12031_ (.A1(_00381_),
    .A2(_02051_),
    .B1(_01956_),
    .B2(_00384_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12032_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02051_),
    .A4(_01956_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12033_ (.A1(_04873_),
    .A2(_04874_),
    .B(_04875_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12034_ (.I(_04876_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12035_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02153_),
    .A4(_02051_),
    .Z(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12036_ (.A1(_04878_),
    .A2(_04744_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12037_ (.A1(_04743_),
    .A2(_04879_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12038_ (.A1(_04877_),
    .A2(_04880_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12039_ (.A1(_00397_),
    .A2(_01693_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12040_ (.A1(_00390_),
    .A2(_01794_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12041_ (.A1(_00393_),
    .A2(_01792_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12042_ (.A1(_04882_),
    .A2(_04883_),
    .A3(_04884_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12043_ (.A1(_04881_),
    .A2(_04885_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12044_ (.A1(_04877_),
    .A2(_04880_),
    .B(_04886_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12045_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02238_),
    .A4(_02236_),
    .Z(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12046_ (.A1(_00378_),
    .A2(_02153_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12047_ (.A1(_00372_),
    .A2(_02238_),
    .B1(_02236_),
    .B2(_00375_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12048_ (.A1(_04888_),
    .A2(_04890_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12049_ (.A1(_04889_),
    .A2(_04891_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12050_ (.A1(_04888_),
    .A2(_04892_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12051_ (.A1(_00369_),
    .A2(_02409_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12052_ (.A1(_00361_),
    .A2(_02584_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12053_ (.A1(_00365_),
    .A2(_02499_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12054_ (.A1(_04895_),
    .A2(_04896_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12055_ (.A1(_04895_),
    .A2(_04896_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12056_ (.A1(_04894_),
    .A2(_04897_),
    .B(_04898_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12057_ (.A1(_04761_),
    .A2(_04763_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12058_ (.A1(_04899_),
    .A2(_04900_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12059_ (.A1(_04899_),
    .A2(_04900_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12060_ (.A1(_04893_),
    .A2(_04901_),
    .B(_04902_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12061_ (.A1(_04753_),
    .A2(_04757_),
    .Z(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12062_ (.A1(_04903_),
    .A2(_04904_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12063_ (.A1(_04903_),
    .A2(_04904_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12064_ (.A1(_04887_),
    .A2(_04905_),
    .B(_04906_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12065_ (.A1(_04755_),
    .A2(_04756_),
    .Z(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12066_ (.A1(_04755_),
    .A2(_04756_),
    .Z(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12067_ (.A1(_04754_),
    .A2(_04908_),
    .B(_04909_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12068_ (.I(_04910_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12069_ (.A1(_04907_),
    .A2(_04911_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12070_ (.A1(_04907_),
    .A2(_04910_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12071_ (.A1(_04887_),
    .A2(_04905_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12072_ (.A1(_04893_),
    .A2(_04901_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12073_ (.A1(_04894_),
    .A2(_04895_),
    .A3(_04896_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12074_ (.A1(_00359_),
    .A2(_02584_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12075_ (.A1(net86),
    .A2(_02762_),
    .B1(_02586_),
    .B2(net83),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12076_ (.A1(net86),
    .A2(net83),
    .A3(_02762_),
    .A4(_02586_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12077_ (.A1(_04917_),
    .A2(_04918_),
    .B(_04919_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12078_ (.A1(_00351_),
    .A2(_02854_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12079_ (.A1(_00354_),
    .A2(_02762_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12080_ (.A1(_04921_),
    .A2(_04922_),
    .A3(_04805_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12081_ (.A1(_04920_),
    .A2(_04923_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12082_ (.A1(_04920_),
    .A2(_04923_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12083_ (.A1(_04916_),
    .A2(_04924_),
    .B(_04925_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12084_ (.A1(_04804_),
    .A2(_04813_),
    .Z(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12085_ (.A1(_04926_),
    .A2(_04927_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12086_ (.A1(_04926_),
    .A2(_04927_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12087_ (.A1(_04915_),
    .A2(_04928_),
    .B(_04929_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12088_ (.A1(_04803_),
    .A2(_04828_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12089_ (.A1(_04930_),
    .A2(_04931_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12090_ (.A1(_04930_),
    .A2(_04931_),
    .Z(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12091_ (.A1(_04914_),
    .A2(_04932_),
    .B(_04933_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12092_ (.A1(_04802_),
    .A2(_04844_),
    .Z(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12093_ (.A1(_04934_),
    .A2(_04935_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12094_ (.A1(_04934_),
    .A2(_04935_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12095_ (.A1(_04913_),
    .A2(_04936_),
    .B(_04937_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12096_ (.A1(_04801_),
    .A2(_04859_),
    .Z(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12097_ (.A1(_04938_),
    .A2(_04939_),
    .Z(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12098_ (.A1(_04938_),
    .A2(_04939_),
    .Z(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12099_ (.A1(_04912_),
    .A2(_04940_),
    .B(_04941_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12100_ (.A1(_04872_),
    .A2(_04942_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12101_ (.A1(_04912_),
    .A2(_04940_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12102_ (.A1(_00387_),
    .A2(_01792_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12103_ (.A1(_00381_),
    .A2(_01956_),
    .B1(_01794_),
    .B2(_00384_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12104_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_01956_),
    .A4(_01794_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12105_ (.A1(_04945_),
    .A2(_04946_),
    .B(_04947_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12106_ (.I(_04948_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12107_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_02051_),
    .A4(_01956_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12108_ (.A1(_04950_),
    .A2(_04874_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12109_ (.A1(_04873_),
    .A2(_04951_),
    .Z(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12110_ (.A1(_04949_),
    .A2(_04952_),
    .Z(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12111_ (.A1(_00397_),
    .A2(_01610_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12112_ (.A1(_00390_),
    .A2(_01792_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12113_ (.A1(_00393_),
    .A2(_01693_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12114_ (.A1(_04954_),
    .A2(_04955_),
    .A3(_04956_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12115_ (.A1(_04953_),
    .A2(_04957_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12116_ (.A1(_04949_),
    .A2(_04952_),
    .B(_04958_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12117_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02236_),
    .A4(_02153_),
    .Z(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12118_ (.A1(_00378_),
    .A2(_02051_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12119_ (.A1(_00372_),
    .A2(_02236_),
    .B1(_02153_),
    .B2(_00375_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12120_ (.A1(_04960_),
    .A2(_04962_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12121_ (.A1(_04961_),
    .A2(_04963_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12122_ (.A1(_04960_),
    .A2(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12123_ (.A1(_00369_),
    .A2(_02238_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12124_ (.A1(_00361_),
    .A2(_02499_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12125_ (.A1(_00365_),
    .A2(_02409_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12126_ (.A1(_04967_),
    .A2(_04968_),
    .Z(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12127_ (.A1(_04967_),
    .A2(_04968_),
    .Z(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12128_ (.A1(_04966_),
    .A2(_04969_),
    .B(_04970_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12129_ (.A1(_04889_),
    .A2(_04891_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12130_ (.A1(_04971_),
    .A2(_04972_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12131_ (.A1(_04971_),
    .A2(_04972_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12132_ (.A1(_04965_),
    .A2(_04973_),
    .B(_04974_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12133_ (.A1(_04881_),
    .A2(_04885_),
    .Z(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12134_ (.A1(_04975_),
    .A2(_04976_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12135_ (.A1(_04975_),
    .A2(_04976_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12136_ (.A1(_04959_),
    .A2(_04977_),
    .B(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12137_ (.A1(_04883_),
    .A2(_04884_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12138_ (.A1(_04883_),
    .A2(_04884_),
    .Z(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12139_ (.A1(_04882_),
    .A2(_04980_),
    .B(_04981_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12140_ (.I(_04982_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12141_ (.A1(_04979_),
    .A2(_04983_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12142_ (.I(_04984_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12143_ (.A1(_04979_),
    .A2(_04982_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12144_ (.A1(_04959_),
    .A2(_04977_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12145_ (.A1(_04965_),
    .A2(_04973_),
    .Z(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12146_ (.A1(_04966_),
    .A2(_04967_),
    .A3(_04968_),
    .Z(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12147_ (.A1(_00359_),
    .A2(_02499_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12148_ (.A1(net66),
    .A2(_02586_),
    .B1(net135),
    .B2(net54),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12149_ (.A1(net66),
    .A2(net54),
    .A3(_02586_),
    .A4(net135),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12150_ (.A1(_04990_),
    .A2(_04991_),
    .B(_04992_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12151_ (.A1(_00351_),
    .A2(_02762_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12152_ (.A1(_00354_),
    .A2(_02586_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12153_ (.A1(_04994_),
    .A2(_04995_),
    .A3(_04917_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12154_ (.A1(_04993_),
    .A2(_04996_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12155_ (.A1(_04993_),
    .A2(_04996_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12156_ (.A1(_04989_),
    .A2(_04997_),
    .B(_04998_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12157_ (.A1(_04916_),
    .A2(_04924_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12158_ (.A1(_04999_),
    .A2(_05000_),
    .Z(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12159_ (.A1(_04999_),
    .A2(_05000_),
    .Z(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12160_ (.A1(_04988_),
    .A2(_05001_),
    .B(_05002_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12161_ (.A1(_04915_),
    .A2(_04928_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12162_ (.A1(_05003_),
    .A2(_05004_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12163_ (.A1(_05003_),
    .A2(_05004_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12164_ (.A1(_04987_),
    .A2(_05005_),
    .B(_05006_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12165_ (.A1(_04914_),
    .A2(_04932_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12166_ (.A1(_05007_),
    .A2(_05008_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12167_ (.A1(_05007_),
    .A2(_05008_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12168_ (.A1(_04986_),
    .A2(_05009_),
    .B(_05010_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12169_ (.A1(_04934_),
    .A2(_04935_),
    .A3(_04913_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12170_ (.A1(_05011_),
    .A2(_05012_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12171_ (.A1(_05011_),
    .A2(_05012_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12172_ (.A1(_04985_),
    .A2(_05013_),
    .B(_05014_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12173_ (.A1(_04944_),
    .A2(_05015_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _12174_ (.A1(_04943_),
    .A2(_05016_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12175_ (.A1(_04397_),
    .A2(_04398_),
    .Z(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12176_ (.A1(_04397_),
    .A2(_04398_),
    .Z(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12177_ (.A1(_04399_),
    .A2(_05018_),
    .B(_05019_),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12178_ (.A1(_00387_),
    .A2(_01693_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12179_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_01794_),
    .A4(_01792_),
    .Z(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12180_ (.A1(_00381_),
    .A2(_01794_),
    .B1(_01792_),
    .B2(_00384_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12181_ (.A1(_05022_),
    .A2(_05023_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12182_ (.A1(_05021_),
    .A2(_05024_),
    .Z(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12183_ (.A1(_05020_),
    .A2(_05025_),
    .Z(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12184_ (.A1(_00397_),
    .A2(_01430_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12185_ (.A1(_00393_),
    .A2(_01524_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12186_ (.A1(_00390_),
    .A2(_01610_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12187_ (.A1(_05027_),
    .A2(_05028_),
    .A3(_05029_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12188_ (.I(_05030_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12189_ (.I(_05025_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12190_ (.A1(_05020_),
    .A2(_05032_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12191_ (.A1(_05026_),
    .A2(_05031_),
    .B(_05033_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12192_ (.A1(_04379_),
    .A2(_04380_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12193_ (.A1(_04379_),
    .A2(_04380_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12194_ (.A1(_04382_),
    .A2(_05035_),
    .B(_05036_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12195_ (.A1(_04367_),
    .A2(_04368_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12196_ (.A1(_04367_),
    .A2(_04368_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12197_ (.A1(_04366_),
    .A2(_05038_),
    .B(_05039_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12198_ (.A1(_00378_),
    .A2(_01956_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12199_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_02153_),
    .A4(_02051_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12200_ (.A1(_00372_),
    .A2(_02153_),
    .B1(_02051_),
    .B2(_00375_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12201_ (.A1(_05042_),
    .A2(_05043_),
    .Z(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12202_ (.A1(_05041_),
    .A2(_05044_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12203_ (.A1(_05040_),
    .A2(_05045_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12204_ (.A1(_05040_),
    .A2(_05045_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12205_ (.A1(_05037_),
    .A2(_05046_),
    .B(_05047_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12206_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_01794_),
    .A4(_01792_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12207_ (.A1(_05021_),
    .A2(_05023_),
    .B(_05049_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12208_ (.I(_05050_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12209_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_01956_),
    .A4(_01794_),
    .Z(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12210_ (.A1(_05052_),
    .A2(_04946_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12211_ (.A1(_04945_),
    .A2(_05053_),
    .Z(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12212_ (.A1(_05051_),
    .A2(_05054_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12213_ (.A1(_00397_),
    .A2(_01524_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12214_ (.A1(_00390_),
    .A2(_01693_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12215_ (.A1(_00393_),
    .A2(_01610_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12216_ (.A1(_05056_),
    .A2(_05057_),
    .A3(_05058_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12217_ (.A1(_05055_),
    .A2(_05059_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12218_ (.A1(_05048_),
    .A2(_05060_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12219_ (.A1(_05048_),
    .A2(_05060_),
    .Z(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12220_ (.A1(_05034_),
    .A2(_05061_),
    .B(_05062_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12221_ (.A1(_05057_),
    .A2(_05058_),
    .Z(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12222_ (.A1(_05057_),
    .A2(_05058_),
    .Z(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12223_ (.A1(_05056_),
    .A2(_05064_),
    .B(_05065_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12224_ (.I(_05066_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12225_ (.A1(_05063_),
    .A2(_05067_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12226_ (.A1(_05063_),
    .A2(_05066_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12227_ (.A1(_04360_),
    .A2(_04364_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12228_ (.A1(_04365_),
    .A2(_04369_),
    .B(_05070_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12229_ (.A1(net87),
    .A2(_02584_),
    .B1(_02499_),
    .B2(net84),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12230_ (.A1(net87),
    .A2(net84),
    .A3(_02584_),
    .A4(_02499_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12231_ (.A1(_04363_),
    .A2(_05072_),
    .B(_05073_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12232_ (.A1(_00354_),
    .A2(_02584_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12233_ (.A1(_00351_),
    .A2(_02586_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12234_ (.A1(_05075_),
    .A2(_05076_),
    .A3(_04990_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12235_ (.A1(_05077_),
    .A2(_05074_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12236_ (.A1(_00369_),
    .A2(_02236_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12237_ (.A1(_00365_),
    .A2(_02238_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12238_ (.A1(_00361_),
    .A2(_02409_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12239_ (.A1(_05079_),
    .A2(_05080_),
    .A3(_05081_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12240_ (.A1(_05078_),
    .A2(_05082_),
    .Z(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12241_ (.A1(_05083_),
    .A2(_05071_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12242_ (.A1(_05037_),
    .A2(_05046_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12243_ (.A1(_05071_),
    .A2(net80),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12244_ (.A1(_05084_),
    .A2(_05085_),
    .B(_05086_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12245_ (.A1(_05074_),
    .A2(_05077_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12246_ (.A1(_05078_),
    .A2(_05082_),
    .B(_05088_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12247_ (.A1(_04989_),
    .A2(_04997_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12248_ (.A1(_05089_),
    .A2(_05090_),
    .Z(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12249_ (.A1(_05041_),
    .A2(_05044_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12250_ (.A1(_05042_),
    .A2(_05092_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12251_ (.A1(_05080_),
    .A2(_05081_),
    .Z(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12252_ (.A1(_05080_),
    .A2(_05081_),
    .Z(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12253_ (.A1(_05079_),
    .A2(_05094_),
    .B(_05095_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12254_ (.A1(_04961_),
    .A2(_04963_),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12255_ (.A1(_05096_),
    .A2(_05097_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12256_ (.A1(_05093_),
    .A2(_05098_),
    .Z(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12257_ (.A1(_05091_),
    .A2(_05099_),
    .Z(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12258_ (.A1(_05087_),
    .A2(_05100_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12259_ (.A1(_05034_),
    .A2(_05061_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12260_ (.A1(_05087_),
    .A2(_05100_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12261_ (.A1(_05101_),
    .A2(_05102_),
    .B(_05103_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12262_ (.A1(_05089_),
    .A2(_05090_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12263_ (.A1(_05091_),
    .A2(_05099_),
    .B(_05105_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12264_ (.A1(_04988_),
    .A2(_05001_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12265_ (.A1(_05106_),
    .A2(_05107_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12266_ (.A1(_05055_),
    .A2(_05059_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12267_ (.A1(_05051_),
    .A2(_05054_),
    .B(_05109_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12268_ (.A1(_05096_),
    .A2(_05097_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12269_ (.A1(_05093_),
    .A2(_05098_),
    .B(_05111_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12270_ (.A1(_04953_),
    .A2(_04957_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12271_ (.A1(_05112_),
    .A2(_05113_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12272_ (.A1(_05110_),
    .A2(_05114_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12273_ (.A1(_05108_),
    .A2(_05115_),
    .Z(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12274_ (.A1(_05104_),
    .A2(_05116_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12275_ (.A1(_05104_),
    .A2(_05116_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12276_ (.A1(_05069_),
    .A2(_05117_),
    .B(_05118_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12277_ (.A1(_05106_),
    .A2(_05107_),
    .Z(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12278_ (.A1(_05108_),
    .A2(_05115_),
    .B(_05120_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12279_ (.A1(_04987_),
    .A2(_05005_),
    .Z(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12280_ (.A1(_05112_),
    .A2(_05113_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12281_ (.A1(_05110_),
    .A2(_05114_),
    .B(_05123_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12282_ (.A1(_04955_),
    .A2(_04956_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12283_ (.A1(_04955_),
    .A2(_04956_),
    .Z(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12284_ (.A1(_04954_),
    .A2(_05125_),
    .B(_05126_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12285_ (.A1(_05124_),
    .A2(_05127_),
    .Z(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12286_ (.A1(_05121_),
    .A2(_05122_),
    .A3(_05128_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12287_ (.A1(_05068_),
    .A2(_05119_),
    .A3(_05129_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12288_ (.I(_04400_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12289_ (.A1(_04396_),
    .A2(_05131_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12290_ (.A1(_04401_),
    .A2(_04406_),
    .B(_05132_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12291_ (.A1(_04378_),
    .A2(_04383_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12292_ (.A1(_04375_),
    .A2(_04384_),
    .B(_05134_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12293_ (.A1(_05026_),
    .A2(_05031_),
    .Z(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12294_ (.A1(_05135_),
    .A2(_05136_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12295_ (.A1(_05135_),
    .A2(_05136_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12296_ (.A1(net94),
    .A2(_05137_),
    .B(_05138_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12297_ (.A1(_05028_),
    .A2(_05029_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12298_ (.A1(_05028_),
    .A2(_05029_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12299_ (.A1(_05027_),
    .A2(_05141_),
    .B(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _12300_ (.I(_05143_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12301_ (.A1(_05140_),
    .A2(_05144_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12302_ (.I(_05145_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12303_ (.A1(_04357_),
    .A2(_04370_),
    .Z(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12304_ (.A1(_04371_),
    .A2(_04385_),
    .B(_05147_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12305_ (.A1(_05084_),
    .A2(_05085_),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12306_ (.A1(_05148_),
    .A2(_05149_),
    .Z(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12307_ (.A1(_05133_),
    .A2(_05135_),
    .A3(_05136_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12308_ (.A1(_04371_),
    .A2(_04385_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12309_ (.A1(_05147_),
    .A2(_05152_),
    .B(net65),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12310_ (.A1(_05150_),
    .A2(_05151_),
    .B(_05153_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12311_ (.A1(_05101_),
    .A2(_05102_),
    .Z(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12312_ (.A1(_05154_),
    .A2(_05155_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12313_ (.A1(_05154_),
    .A2(_05155_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12314_ (.A1(_05146_),
    .A2(_05156_),
    .B(_05157_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12315_ (.A1(_05069_),
    .A2(_05117_),
    .Z(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12316_ (.A1(_05158_),
    .A2(_05159_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12317_ (.A1(_05158_),
    .A2(_05159_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _12318_ (.A1(_05140_),
    .A2(_05144_),
    .A3(_05161_),
    .B(_05162_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12319_ (.A1(_05130_),
    .A2(_05163_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12320_ (.A1(_05140_),
    .A2(_05144_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12321_ (.A1(_05158_),
    .A2(_05159_),
    .Z(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12322_ (.A1(_05165_),
    .A2(_05166_),
    .Z(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12323_ (.A1(_04393_),
    .A2(_04407_),
    .Z(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12324_ (.A1(_04393_),
    .A2(_04407_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12325_ (.A1(_04391_),
    .A2(_05168_),
    .B(_05169_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12326_ (.A1(_00397_),
    .A2(_01249_),
    .A3(_04405_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12327_ (.A1(_04403_),
    .A2(_04404_),
    .B(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12328_ (.I(_05173_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12329_ (.A1(_05170_),
    .A2(_05174_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _12330_ (.I(_05175_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12331_ (.A1(_05170_),
    .A2(_05174_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12332_ (.A1(_05176_),
    .A2(_05177_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12333_ (.A1(_04371_),
    .A2(_04385_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _12334_ (.A1(_05152_),
    .A2(_04387_),
    .A3(_05179_),
    .B1(_04388_),
    .B2(_04408_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12335_ (.A1(_05151_),
    .A2(_05150_),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12336_ (.A1(_05180_),
    .A2(_05181_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12337_ (.A1(_05180_),
    .A2(_05181_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12338_ (.A1(_05178_),
    .A2(_05183_),
    .B(_05184_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12339_ (.A1(_05154_),
    .A2(_05155_),
    .A3(_05145_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12340_ (.A1(_05185_),
    .A2(_05186_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12341_ (.A1(_05185_),
    .A2(_05186_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12342_ (.A1(_05176_),
    .A2(_05187_),
    .B(_05188_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12343_ (.A1(_05167_),
    .A2(_05189_),
    .Z(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12344_ (.A1(_05164_),
    .A2(_05190_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12345_ (.A1(_05176_),
    .A2(_05185_),
    .A3(_05186_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12346_ (.A1(_04348_),
    .A2(_04351_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12347_ (.I(_04352_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12348_ (.A1(_04355_),
    .A2(_04409_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12349_ (.A1(_05195_),
    .A2(_04410_),
    .B(_05196_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12350_ (.A1(_05180_),
    .A2(_05181_),
    .A3(_05178_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12351_ (.A1(_05198_),
    .A2(_05197_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12352_ (.A1(_05197_),
    .A2(_05198_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12353_ (.A1(_05194_),
    .A2(net82),
    .B(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12354_ (.A1(_05192_),
    .A2(_05201_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12355_ (.A1(_05192_),
    .A2(_05201_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12356_ (.A1(_05194_),
    .A2(_05199_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12357_ (.A1(_04345_),
    .A2(_04411_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12358_ (.A1(_04224_),
    .A2(_04412_),
    .B(_05206_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12359_ (.A1(_05205_),
    .A2(_05207_),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _12360_ (.A1(_05202_),
    .A2(_05203_),
    .A3(_05208_),
    .Z(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12361_ (.A1(_05011_),
    .A2(_05012_),
    .Z(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12362_ (.A1(_04985_),
    .A2(_05210_),
    .Z(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12363_ (.I(_05127_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12364_ (.A1(_05124_),
    .A2(_05212_),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12365_ (.A1(_05121_),
    .A2(_05122_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12366_ (.A1(_05121_),
    .A2(_05122_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12367_ (.A1(_05128_),
    .A2(_05214_),
    .B(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12368_ (.A1(_04986_),
    .A2(_05009_),
    .Z(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12369_ (.A1(_05217_),
    .A2(_05218_),
    .Z(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12370_ (.A1(_05217_),
    .A2(_05218_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12371_ (.A1(_05213_),
    .A2(_05219_),
    .B(_05220_),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12372_ (.A1(_05211_),
    .A2(_05221_),
    .Z(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12373_ (.A1(_05213_),
    .A2(_05219_),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12374_ (.A1(_05119_),
    .A2(_05129_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12375_ (.A1(_05119_),
    .A2(_05129_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _12376_ (.A1(_05063_),
    .A2(_05067_),
    .A3(_05224_),
    .B(_05225_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12377_ (.A1(_05223_),
    .A2(_05227_),
    .Z(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _12378_ (.A1(_05222_),
    .A2(_05228_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _12379_ (.A1(_05017_),
    .A2(_05191_),
    .A3(_05209_),
    .A4(_05229_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12380_ (.A1(_05211_),
    .A2(_05221_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12381_ (.A1(_05223_),
    .A2(_05227_),
    .Z(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12382_ (.A1(_05211_),
    .A2(_05221_),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12383_ (.A1(_05231_),
    .A2(_05232_),
    .B(_05233_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12384_ (.A1(_04872_),
    .A2(_04942_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12385_ (.A1(_04984_),
    .A2(_05210_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12386_ (.A1(_05014_),
    .A2(_05236_),
    .B(_04944_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12387_ (.A1(_04872_),
    .A2(_04942_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12388_ (.A1(_05235_),
    .A2(_05238_),
    .B(_05239_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12389_ (.A1(_05017_),
    .A2(_05234_),
    .B(_05240_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12390_ (.A1(_05192_),
    .A2(_05201_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _12391_ (.A1(_05192_),
    .A2(_05201_),
    .B1(_05205_),
    .B2(_05207_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12392_ (.A1(_05164_),
    .A2(_05190_),
    .A3(_05242_),
    .A4(_05243_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12393_ (.A1(_05130_),
    .A2(_05163_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _12394_ (.A1(_05130_),
    .A2(_05163_),
    .B(_05167_),
    .C(_05189_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12395_ (.A1(_05245_),
    .A2(_05246_),
    .Z(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _12396_ (.A1(_05244_),
    .A2(_05247_),
    .B(_05229_),
    .C(_05017_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _12397_ (.A1(_04742_),
    .A2(_05230_),
    .B(_05241_),
    .C(_05249_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12398_ (.I(_04869_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12399_ (.A1(_04863_),
    .A2(_04864_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12400_ (.A1(_04863_),
    .A2(_04864_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12401_ (.A1(_04870_),
    .A2(_05252_),
    .B(_05253_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12402_ (.A1(_04168_),
    .A2(_04146_),
    .Z(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12403_ (.A1(_05254_),
    .A2(_05255_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12404_ (.A1(_05254_),
    .A2(_05255_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _12405_ (.A1(_04866_),
    .A2(_05251_),
    .A3(_05256_),
    .B(_05257_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12406_ (.A1(_04141_),
    .A2(_04145_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12407_ (.A1(_05259_),
    .A2(_04172_),
    .Z(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12408_ (.A1(_05258_),
    .A2(_05260_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12409_ (.A1(_04866_),
    .A2(_05251_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12410_ (.A1(_05254_),
    .A2(_05255_),
    .Z(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12411_ (.A1(_05262_),
    .A2(_05263_),
    .Z(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12412_ (.A1(_04861_),
    .A2(_04871_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12413_ (.A1(_04861_),
    .A2(_04871_),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12414_ (.A1(_04800_),
    .A2(_05265_),
    .B(_05266_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12415_ (.A1(_05264_),
    .A2(_05267_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12416_ (.A1(_05261_),
    .A2(_05268_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12417_ (.A1(_05262_),
    .A2(_05263_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12418_ (.A1(_05257_),
    .A2(_05271_),
    .B(_05260_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12419_ (.A1(_05264_),
    .A2(_05267_),
    .Z(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12420_ (.A1(_05257_),
    .A2(_05271_),
    .A3(_05260_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12421_ (.A1(_05272_),
    .A2(_05273_),
    .B(_05274_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12422_ (.A1(_05250_),
    .A2(_05270_),
    .B(_05275_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12423_ (.A1(_04106_),
    .A2(_04173_),
    .Z(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12424_ (.A1(_04174_),
    .A2(_05276_),
    .B(_05277_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12425_ (.A1(_04105_),
    .A2(_05278_),
    .Z(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12426_ (.A1(_04174_),
    .A2(_05276_),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _12427_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-15] ),
    .A2(_05281_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12428_ (.A1(_05223_),
    .A2(_05227_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12429_ (.A1(_05191_),
    .A2(_05209_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _12430_ (.A1(_05164_),
    .A2(_05190_),
    .A3(_05242_),
    .A4(_05243_),
    .Z(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12431_ (.A1(_05245_),
    .A2(_05246_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _12432_ (.A1(_04742_),
    .A2(_05284_),
    .B(_05285_),
    .C(_05286_),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12433_ (.A1(_05223_),
    .A2(_05227_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12434_ (.A1(_05283_),
    .A2(_05287_),
    .B(_05288_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12435_ (.A1(_05222_),
    .A2(_05289_),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12436_ (.A1(_05283_),
    .A2(_05287_),
    .Z(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12437_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-20] ),
    .A2(_05290_),
    .B1(_05292_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-21] ),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12438_ (.A1(_05242_),
    .A2(_05243_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _12439_ (.A1(_04740_),
    .A2(_04741_),
    .A3(_05209_),
    .B(_05294_),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12440_ (.A1(_05190_),
    .A2(_05295_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12441_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-23] ),
    .A2(_05296_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _12442_ (.A1(_04740_),
    .A2(_04741_),
    .Z(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _12443_ (.A1(_04740_),
    .A2(_04741_),
    .A3(_05208_),
    .B(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-25] ),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12444_ (.A1(_05298_),
    .A2(_05208_),
    .B(_05299_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12445_ (.A1(_05202_),
    .A2(_05203_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _12446_ (.A1(_04740_),
    .A2(_04741_),
    .A3(_05208_),
    .B1(_05207_),
    .B2(_05205_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12447_ (.A1(_05301_),
    .A2(_05303_),
    .Z(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12448_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-24] ),
    .A2(_05300_),
    .B(_05304_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12449_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-24] ),
    .A2(_05300_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _12450_ (.A1(_05297_),
    .A2(_05305_),
    .A3(_05306_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12451_ (.A1(_05167_),
    .A2(_05189_),
    .Z(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12452_ (.A1(_05190_),
    .A2(_05295_),
    .B(_05308_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12453_ (.A1(_05164_),
    .A2(_05309_),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12454_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-23] ),
    .A2(_05296_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12455_ (.A1(_03763_),
    .A2(_05310_),
    .B(_05311_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12456_ (.A1(_03763_),
    .A2(_05310_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _12457_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-21] ),
    .A2(_05292_),
    .B1(_05307_),
    .B2(_05312_),
    .C(_05314_),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12458_ (.A1(_05287_),
    .A2(_05229_),
    .B(_05234_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12459_ (.A1(_05016_),
    .A2(_05316_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _12460_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-19] ),
    .A2(_05317_),
    .B1(_05290_),
    .B2(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-20] ),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12461_ (.A1(_05293_),
    .A2(_05315_),
    .B(_05318_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12462_ (.A1(_05016_),
    .A2(_05316_),
    .B(_05238_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12463_ (.A1(_04943_),
    .A2(_05320_),
    .Z(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12464_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-19] ),
    .A2(_05317_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12465_ (.A1(_03768_),
    .A2(_05321_),
    .B(_05322_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12466_ (.A1(_03768_),
    .A2(_05321_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _12467_ (.A1(_05319_),
    .A2(_05323_),
    .B(_05325_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _12468_ (.A1(_05017_),
    .A2(_05191_),
    .A3(_05209_),
    .A4(_05229_),
    .Z(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12469_ (.A1(_04943_),
    .A2(_05016_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12470_ (.A1(_05211_),
    .A2(_05221_),
    .Z(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12471_ (.A1(_05211_),
    .A2(_05221_),
    .Z(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12472_ (.A1(_05329_),
    .A2(_05288_),
    .B(_05330_),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _12473_ (.A1(_05235_),
    .A2(_05238_),
    .B1(_05328_),
    .B2(_05331_),
    .C(_05239_),
    .ZN(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12474_ (.A1(_05222_),
    .A2(_05228_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _12475_ (.A1(_05285_),
    .A2(_05286_),
    .B(_05333_),
    .C(_05328_),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _12476_ (.A1(_05298_),
    .A2(_05327_),
    .B(_05332_),
    .C(_05334_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12477_ (.A1(_05336_),
    .A2(_05268_),
    .B(_05273_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12478_ (.A1(_05261_),
    .A2(_05337_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12479_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-16] ),
    .A2(_05338_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12480_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-16] ),
    .A2(_05338_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12481_ (.A1(_05336_),
    .A2(_05268_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12482_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-17] ),
    .A2(_05341_),
    .Z(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12483_ (.I(_05342_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12484_ (.A1(_05343_),
    .A2(_05340_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12485_ (.A1(_05339_),
    .A2(_05344_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12486_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-17] ),
    .A2(_05341_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12487_ (.A1(_05339_),
    .A2(_05347_),
    .B(_05340_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12488_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-15] ),
    .A2(_05281_),
    .B(_05348_),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12489_ (.A1(_05326_),
    .A2(_05345_),
    .B(_05349_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12490_ (.A1(_05282_),
    .A2(_05350_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12491_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-14] ),
    .A2(_05279_),
    .A3(_05351_),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12492_ (.I0(net20),
    .I1(_05352_),
    .S(_05171_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12493_ (.I(_05353_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12494_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-15] ),
    .A2(_05281_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12495_ (.A1(_03773_),
    .A2(_05279_),
    .B(_05354_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12496_ (.A1(_03773_),
    .A2(_05279_),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12497_ (.A1(_05356_),
    .A2(_05282_),
    .A3(_05339_),
    .A4(_05344_),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12498_ (.A1(_05282_),
    .A2(_05348_),
    .B(_05355_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12499_ (.I(_05356_),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _12500_ (.A1(_05326_),
    .A2(_05355_),
    .A3(_05357_),
    .B1(_05358_),
    .B2(_05359_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12501_ (.A1(_03981_),
    .A2(_04033_),
    .Z(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12502_ (.A1(_03979_),
    .A2(_04034_),
    .B(_05361_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12503_ (.A1(_04017_),
    .A2(_04031_),
    .Z(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12504_ (.A1(_04017_),
    .A2(_04031_),
    .Z(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12505_ (.A1(_04015_),
    .A2(_05363_),
    .B(_05364_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12506_ (.A1(_00397_),
    .A2(_02409_),
    .A3(_04021_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12507_ (.A1(_04019_),
    .A2(_04020_),
    .B(_05367_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12508_ (.A1(_05365_),
    .A2(_05368_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12509_ (.A1(_03930_),
    .A2(_03946_),
    .Z(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12510_ (.A1(_03982_),
    .A2(_05370_),
    .B(_04011_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12511_ (.A1(_04012_),
    .A2(_04032_),
    .B(_05371_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12512_ (.A1(_03985_),
    .A2(_03998_),
    .Z(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12513_ (.A1(_03999_),
    .A2(_04010_),
    .B(_05373_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12514_ (.A1(_03988_),
    .A2(_03992_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12515_ (.A1(_03993_),
    .A2(_03997_),
    .B(_05375_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12516_ (.A1(_03556_),
    .A2(net86),
    .B1(net83),
    .B2(_03485_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12517_ (.A1(_03556_),
    .A2(net86),
    .A3(net83),
    .A4(_03485_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12518_ (.A1(_03989_),
    .A2(_05377_),
    .B(_05378_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12519_ (.A1(_03485_),
    .A2(_00359_),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12520_ (.A1(_03556_),
    .A2(_00354_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12521_ (.A1(net86),
    .A2(_03558_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12522_ (.A1(_05380_),
    .A2(_05381_),
    .A3(_05382_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12523_ (.A1(_05379_),
    .A2(_05383_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12524_ (.A1(_03266_),
    .A2(_00369_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12525_ (.A1(_03340_),
    .A2(_00365_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12526_ (.A1(net148),
    .A2(_00361_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12527_ (.A1(_05385_),
    .A2(_05386_),
    .A3(_05388_),
    .Z(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12528_ (.A1(_05384_),
    .A2(_05389_),
    .Z(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12529_ (.A1(_05376_),
    .A2(_05390_),
    .Z(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12530_ (.A1(_04006_),
    .A2(_04007_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12531_ (.A1(_04006_),
    .A2(_04007_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12532_ (.A1(_04005_),
    .A2(_05392_),
    .B(_05393_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12533_ (.A1(_03995_),
    .A2(_03996_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12534_ (.A1(_03995_),
    .A2(_03996_),
    .Z(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12535_ (.A1(_03994_),
    .A2(_05395_),
    .B(_05396_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12536_ (.A1(_02940_),
    .A2(_00378_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12537_ (.A1(_03018_),
    .A2(_00375_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12538_ (.A1(_03189_),
    .A2(_00372_),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12539_ (.A1(_05399_),
    .A2(_05400_),
    .A3(_05401_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12540_ (.A1(_05397_),
    .A2(_05402_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12541_ (.A1(_05394_),
    .A2(_05403_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12542_ (.A1(_05374_),
    .A2(_05391_),
    .A3(_05404_),
    .Z(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12543_ (.I(_04029_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12544_ (.A1(_04025_),
    .A2(_05406_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12545_ (.A1(_04022_),
    .A2(_04030_),
    .B(_05407_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12546_ (.A1(_04003_),
    .A2(_04008_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12547_ (.A1(_04000_),
    .A2(_04009_),
    .B(_05410_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12548_ (.A1(_02499_),
    .A2(_00397_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12549_ (.A1(net135),
    .A2(_00393_),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12550_ (.A1(_02586_),
    .A2(_00390_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12551_ (.A1(_05413_),
    .A2(_05414_),
    .Z(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12552_ (.A1(_05412_),
    .A2(_05415_),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12553_ (.A1(_04027_),
    .A2(_04028_),
    .Z(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12554_ (.A1(_04027_),
    .A2(_04028_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12555_ (.A1(_04026_),
    .A2(_05417_),
    .B(_05418_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12556_ (.A1(_02762_),
    .A2(_00387_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12557_ (.A1(_02854_),
    .A2(_00384_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12558_ (.A1(_02938_),
    .A2(_00381_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12559_ (.A1(_05421_),
    .A2(_05422_),
    .A3(_05423_),
    .Z(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12560_ (.A1(_05419_),
    .A2(_05424_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12561_ (.A1(_05416_),
    .A2(_05425_),
    .Z(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12562_ (.A1(_05411_),
    .A2(_05426_),
    .Z(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12563_ (.A1(_05408_),
    .A2(_05427_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12564_ (.A1(_05428_),
    .A2(_05405_),
    .Z(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12565_ (.A1(_05372_),
    .A2(_05429_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12566_ (.A1(_05430_),
    .A2(_05369_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12567_ (.A1(_05362_),
    .A2(_05432_),
    .Z(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12568_ (.A1(_03977_),
    .A2(_05433_),
    .Z(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12569_ (.A1(_03971_),
    .A2(_04035_),
    .Z(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12570_ (.A1(_03971_),
    .A2(_04035_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12571_ (.A1(_03850_),
    .A2(_05435_),
    .B(_05436_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12572_ (.A1(_05434_),
    .A2(_05437_),
    .Z(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12573_ (.A1(_04105_),
    .A2(_04174_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12574_ (.A1(_04036_),
    .A2(_04104_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12575_ (.A1(_05440_),
    .A2(_05277_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _12576_ (.A1(_04036_),
    .A2(_04104_),
    .B1(_05275_),
    .B2(_05439_),
    .C(_05441_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12577_ (.I(_05443_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _12578_ (.A1(_05250_),
    .A2(_05270_),
    .A3(_05439_),
    .B(_05444_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12579_ (.A1(_05438_),
    .A2(net145),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12580_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-13] ),
    .A2(_05446_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12581_ (.A1(_05360_),
    .A2(_05447_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12582_ (.A1(_05360_),
    .A2(_05447_),
    .B(_05182_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12583_ (.A1(_05280_),
    .A2(net27),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12584_ (.A1(_05448_),
    .A2(_05449_),
    .B(_05450_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12585_ (.I(_05365_),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12586_ (.A1(_05451_),
    .A2(_05368_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12587_ (.A1(_05372_),
    .A2(_05429_),
    .ZN(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12588_ (.A1(_05369_),
    .A2(_05430_),
    .B(_05454_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12589_ (.A1(_05411_),
    .A2(_05426_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12590_ (.A1(_05408_),
    .A2(_05427_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12591_ (.A1(_05456_),
    .A2(_05457_),
    .ZN(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12592_ (.A1(_02499_),
    .A2(_00397_),
    .A3(_05415_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12593_ (.A1(_05413_),
    .A2(_05414_),
    .B(_05459_),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12594_ (.A1(_05458_),
    .A2(_05460_),
    .Z(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12595_ (.A1(_05391_),
    .A2(_05404_),
    .Z(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12596_ (.A1(_05391_),
    .A2(_05404_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _12597_ (.A1(net93),
    .A2(_05462_),
    .A3(_05464_),
    .B1(_05405_),
    .B2(_05428_),
    .ZN(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12598_ (.A1(_05376_),
    .A2(_05390_),
    .Z(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12599_ (.A1(_05391_),
    .A2(_05404_),
    .B(_05466_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12600_ (.A1(_05379_),
    .A2(_05383_),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12601_ (.A1(_05384_),
    .A2(_05389_),
    .B(_05468_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12602_ (.A1(_03556_),
    .A2(net54),
    .B1(_03558_),
    .B2(net66),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12603_ (.A1(_03556_),
    .A2(net66),
    .A3(net54),
    .A4(_03558_),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12604_ (.A1(_05380_),
    .A2(_05470_),
    .B(_05471_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12605_ (.A1(_03556_),
    .A2(_00359_),
    .ZN(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12606_ (.A1(net84),
    .A2(_03558_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12607_ (.A1(net66),
    .A2(_03679_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12608_ (.A1(_05473_),
    .A2(_05475_),
    .A3(_05476_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12609_ (.A1(_05472_),
    .A2(_05477_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12610_ (.A1(_03340_),
    .A2(_00369_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12611_ (.A1(_03485_),
    .A2(net148),
    .A3(_00361_),
    .A4(_00365_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12612_ (.A1(_03485_),
    .A2(_00361_),
    .B1(_00365_),
    .B2(net148),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12613_ (.A1(_05480_),
    .A2(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12614_ (.A1(_05479_),
    .A2(_05482_),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12615_ (.A1(_05478_),
    .A2(_05483_),
    .Z(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12616_ (.A1(_05469_),
    .A2(_05484_),
    .Z(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12617_ (.A1(_05400_),
    .A2(_05401_),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12618_ (.A1(_05400_),
    .A2(_05401_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12619_ (.A1(_05399_),
    .A2(_05487_),
    .B(_05488_),
    .ZN(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12620_ (.A1(_05386_),
    .A2(_05388_),
    .Z(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12621_ (.A1(_05386_),
    .A2(_05388_),
    .Z(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12622_ (.A1(_05385_),
    .A2(_05490_),
    .B(_05491_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12623_ (.A1(_03018_),
    .A2(_00378_),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12624_ (.A1(_03189_),
    .A2(_00375_),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12625_ (.A1(_03266_),
    .A2(_00372_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12626_ (.A1(_05494_),
    .A2(_05495_),
    .Z(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12627_ (.A1(_05493_),
    .A2(_05497_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12628_ (.A1(_05492_),
    .A2(_05498_),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12629_ (.A1(_05489_),
    .A2(_05499_),
    .Z(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12630_ (.A1(_05486_),
    .A2(_05500_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12631_ (.A1(_05467_),
    .A2(_05501_),
    .Z(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12632_ (.I(_05424_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12633_ (.A1(_05419_),
    .A2(_05503_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12634_ (.A1(_05416_),
    .A2(_05425_),
    .B(_05504_),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12635_ (.A1(_05397_),
    .A2(_05402_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12636_ (.A1(_05394_),
    .A2(_05403_),
    .B(_05506_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12637_ (.A1(net135),
    .A2(_00397_),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12638_ (.A1(_02586_),
    .A2(_00393_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12639_ (.A1(_02762_),
    .A2(_00390_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12640_ (.A1(_05510_),
    .A2(_05511_),
    .Z(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12641_ (.A1(_05509_),
    .A2(_05512_),
    .Z(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12642_ (.A1(_05422_),
    .A2(_05423_),
    .Z(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12643_ (.A1(_05422_),
    .A2(_05423_),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12644_ (.A1(_05421_),
    .A2(_05514_),
    .B(_05515_),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12645_ (.A1(_02854_),
    .A2(_00387_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12646_ (.A1(_02938_),
    .A2(_00384_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12647_ (.A1(_02940_),
    .A2(_00381_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12648_ (.A1(_05517_),
    .A2(_05519_),
    .A3(_05520_),
    .Z(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12649_ (.A1(_05516_),
    .A2(_05521_),
    .Z(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12650_ (.A1(_05513_),
    .A2(_05522_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12651_ (.A1(_05505_),
    .A2(_05508_),
    .A3(_05523_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12652_ (.A1(_05502_),
    .A2(_05524_),
    .Z(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12653_ (.A1(_05465_),
    .A2(_05525_),
    .Z(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12654_ (.A1(_05461_),
    .A2(_05526_),
    .Z(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12655_ (.A1(_05453_),
    .A2(_05455_),
    .A3(_05527_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12656_ (.I(_05528_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12657_ (.A1(_05362_),
    .A2(_05432_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12658_ (.A1(_03977_),
    .A2(_05433_),
    .B(_05531_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12659_ (.A1(_05434_),
    .A2(_05437_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12660_ (.A1(_05438_),
    .A2(_05445_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12661_ (.A1(_05533_),
    .A2(_05534_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12662_ (.A1(_05530_),
    .A2(_05532_),
    .A3(_05535_),
    .Z(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12663_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-12] ),
    .A2(_05536_),
    .Z(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12664_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-13] ),
    .A2(_05446_),
    .Z(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12665_ (.A1(_05538_),
    .A2(_05448_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12666_ (.A1(_05537_),
    .A2(_05539_),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12667_ (.A1(_05280_),
    .A2(net28),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12668_ (.A1(_05822_),
    .A2(_05541_),
    .B(_05542_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12669_ (.A1(_05822_),
    .A2(net29),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12670_ (.A1(_05458_),
    .A2(_05460_),
    .Z(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12671_ (.A1(_05465_),
    .A2(_05525_),
    .Z(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12672_ (.A1(_05461_),
    .A2(_05526_),
    .B(_05545_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12673_ (.A1(_05508_),
    .A2(_05523_),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12674_ (.A1(_05508_),
    .A2(_05523_),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12675_ (.A1(_05505_),
    .A2(_05547_),
    .B(_05548_),
    .ZN(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12676_ (.A1(_05510_),
    .A2(_05511_),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12677_ (.A1(net135),
    .A2(_00397_),
    .A3(_05512_),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12678_ (.A1(_05551_),
    .A2(_05552_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12679_ (.A1(_05549_),
    .A2(_05553_),
    .Z(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12680_ (.A1(_05466_),
    .A2(_05462_),
    .B(_05501_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12681_ (.A1(_05502_),
    .A2(_05524_),
    .B(_05555_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12682_ (.A1(_05469_),
    .A2(_05484_),
    .Z(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12683_ (.A1(_05486_),
    .A2(_05500_),
    .B(_05557_),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12684_ (.A1(_05472_),
    .A2(_05477_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12685_ (.A1(_05478_),
    .A2(_05483_),
    .B(_05559_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12686_ (.A1(_00354_),
    .A2(_03558_),
    .B1(_03679_),
    .B2(net87),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12687_ (.A1(net87),
    .A2(_00354_),
    .A3(_03558_),
    .A4(_03679_),
    .ZN(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12688_ (.A1(_05473_),
    .A2(_05562_),
    .B(_05563_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12689_ (.A1(_00359_),
    .A2(_03558_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12690_ (.A1(net86),
    .A2(net84),
    .A3(_03679_),
    .A4(_03725_),
    .Z(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12691_ (.A1(net54),
    .A2(_03679_),
    .B1(_03725_),
    .B2(net86),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12692_ (.A1(_05566_),
    .A2(_05567_),
    .ZN(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12693_ (.A1(_05564_),
    .A2(_05565_),
    .A3(_05568_),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12694_ (.A1(net148),
    .A2(_00369_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12695_ (.A1(_03485_),
    .A2(_00365_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12696_ (.A1(_03556_),
    .A2(_00361_),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12697_ (.A1(_05570_),
    .A2(_05571_),
    .A3(_05573_),
    .Z(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12698_ (.A1(_05569_),
    .A2(_05574_),
    .Z(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12699_ (.A1(_05560_),
    .A2(_05575_),
    .Z(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12700_ (.A1(_05494_),
    .A2(_05495_),
    .Z(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12701_ (.A1(_03018_),
    .A2(_00378_),
    .A3(_05497_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12702_ (.A1(_05577_),
    .A2(_05578_),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12703_ (.I(_05480_),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12704_ (.A1(_05479_),
    .A2(_05481_),
    .B(_05580_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12705_ (.A1(_03189_),
    .A2(_00378_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12706_ (.A1(_03266_),
    .A2(_00375_),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12707_ (.A1(_03340_),
    .A2(_00372_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12708_ (.A1(_05584_),
    .A2(_05585_),
    .Z(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12709_ (.A1(_05582_),
    .A2(_05586_),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12710_ (.A1(_05581_),
    .A2(_05587_),
    .Z(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12711_ (.A1(_05579_),
    .A2(_05588_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12712_ (.A1(_05576_),
    .A2(_05589_),
    .Z(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12713_ (.A1(_05558_),
    .A2(_05590_),
    .Z(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12714_ (.I(_05521_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12715_ (.A1(_05516_),
    .A2(_05592_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12716_ (.A1(_05513_),
    .A2(_05522_),
    .B(_05593_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12717_ (.A1(_05492_),
    .A2(_05498_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12718_ (.A1(_05489_),
    .A2(_05499_),
    .B(_05596_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12719_ (.A1(_02586_),
    .A2(_00397_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12720_ (.A1(_02762_),
    .A2(_00393_),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12721_ (.A1(_02854_),
    .A2(_00390_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12722_ (.A1(_05599_),
    .A2(_05600_),
    .Z(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12723_ (.A1(_05598_),
    .A2(_05601_),
    .Z(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12724_ (.A1(_05519_),
    .A2(_05520_),
    .Z(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12725_ (.A1(_05519_),
    .A2(_05520_),
    .Z(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12726_ (.A1(_05517_),
    .A2(_05603_),
    .B(_05604_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12727_ (.A1(_02938_),
    .A2(_00387_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12728_ (.A1(_02940_),
    .A2(_00384_),
    .ZN(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12729_ (.A1(_03018_),
    .A2(_00381_),
    .ZN(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12730_ (.A1(_05607_),
    .A2(_05608_),
    .A3(_05609_),
    .Z(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12731_ (.A1(_05606_),
    .A2(_05610_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12732_ (.A1(_05602_),
    .A2(_05611_),
    .Z(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12733_ (.A1(_05595_),
    .A2(_05597_),
    .A3(_05612_),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12734_ (.A1(_05591_),
    .A2(_05613_),
    .Z(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12735_ (.A1(_05556_),
    .A2(_05614_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12736_ (.A1(_05554_),
    .A2(_05615_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12737_ (.A1(_05546_),
    .A2(_05617_),
    .Z(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12738_ (.A1(_05544_),
    .A2(_05618_),
    .Z(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12739_ (.A1(_05455_),
    .A2(_05527_),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12740_ (.A1(_05455_),
    .A2(_05527_),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12741_ (.A1(_05453_),
    .A2(_05620_),
    .B(_05621_),
    .ZN(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12742_ (.A1(_05619_),
    .A2(_05622_),
    .ZN(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12743_ (.A1(_05530_),
    .A2(_05532_),
    .Z(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12744_ (.A1(_05530_),
    .A2(_05532_),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12745_ (.A1(_05438_),
    .A2(_05624_),
    .A3(_05625_),
    .Z(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12746_ (.A1(_05530_),
    .A2(_05532_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12747_ (.A1(_05533_),
    .A2(_05624_),
    .B(_05628_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12748_ (.A1(_05445_),
    .A2(_05626_),
    .B(_05629_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12749_ (.A1(_05623_),
    .A2(_05630_),
    .Z(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12750_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-11] ),
    .A2(_05631_),
    .ZN(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12751_ (.A1(_05447_),
    .A2(_05537_),
    .Z(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12752_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-12] ),
    .A2(_05536_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12753_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-12] ),
    .A2(_05536_),
    .B(_05538_),
    .ZN(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12754_ (.A1(_05634_),
    .A2(_05635_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12755_ (.A1(_05360_),
    .A2(_05633_),
    .B(_05636_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12756_ (.A1(_05632_),
    .A2(_05637_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12757_ (.A1(_05632_),
    .A2(_05637_),
    .Z(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12758_ (.A1(_05387_),
    .A2(_05638_),
    .A3(_05639_),
    .ZN(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12759_ (.A1(_05543_),
    .A2(_05640_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12760_ (.A1(_05551_),
    .A2(_05552_),
    .B(_05549_),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12761_ (.A1(_05556_),
    .A2(_05614_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12762_ (.A1(_05554_),
    .A2(_05615_),
    .B(_05642_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12763_ (.A1(_05597_),
    .A2(_05612_),
    .Z(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12764_ (.A1(_05597_),
    .A2(_05612_),
    .Z(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12765_ (.A1(_05595_),
    .A2(_05644_),
    .B(_05645_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12766_ (.A1(_05599_),
    .A2(_05600_),
    .Z(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12767_ (.A1(_02586_),
    .A2(_00397_),
    .A3(_05601_),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12768_ (.A1(_05648_),
    .A2(_05649_),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12769_ (.A1(_05646_),
    .A2(_05650_),
    .Z(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12770_ (.I(_05558_),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12771_ (.A1(_05652_),
    .A2(_05590_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12772_ (.A1(_05591_),
    .A2(_05613_),
    .B(_05653_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12773_ (.A1(_05560_),
    .A2(_05575_),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12774_ (.A1(_05576_),
    .A2(_05589_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12775_ (.A1(_05655_),
    .A2(_05656_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12776_ (.I(_05565_),
    .ZN(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12777_ (.A1(_05659_),
    .A2(_05568_),
    .Z(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12778_ (.A1(_05564_),
    .A2(_05660_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12779_ (.A1(_05569_),
    .A2(_05574_),
    .B(_05661_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12780_ (.A1(_05659_),
    .A2(_05568_),
    .B(_05566_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12781_ (.A1(net83),
    .A2(_03725_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12782_ (.A1(net86),
    .A2(_03727_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12783_ (.A1(net70),
    .A2(_03679_),
    .ZN(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12784_ (.A1(_05664_),
    .A2(_05665_),
    .A3(_05666_),
    .Z(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12785_ (.A1(_05663_),
    .A2(_05667_),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12786_ (.A1(_03485_),
    .A2(_00369_),
    .ZN(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12787_ (.A1(_03556_),
    .A2(_00365_),
    .ZN(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12788_ (.A1(_00361_),
    .A2(_03558_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12789_ (.A1(_05670_),
    .A2(_05671_),
    .A3(_05672_),
    .Z(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12790_ (.A1(_05668_),
    .A2(_05673_),
    .Z(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12791_ (.A1(_05662_),
    .A2(_05674_),
    .Z(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12792_ (.A1(_05584_),
    .A2(_05585_),
    .Z(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12793_ (.A1(_03189_),
    .A2(_00378_),
    .A3(_05586_),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12794_ (.A1(_05571_),
    .A2(_05573_),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12795_ (.A1(_05571_),
    .A2(_05573_),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12796_ (.A1(_05570_),
    .A2(_05678_),
    .B(_05679_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12797_ (.A1(_03266_),
    .A2(_00378_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12798_ (.A1(_03340_),
    .A2(_00375_),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12799_ (.A1(net147),
    .A2(_00372_),
    .ZN(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12800_ (.A1(_05682_),
    .A2(_05683_),
    .A3(_05684_),
    .Z(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12801_ (.A1(_05681_),
    .A2(_05685_),
    .Z(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12802_ (.A1(_05676_),
    .A2(_05677_),
    .B(_05686_),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12803_ (.A1(_05676_),
    .A2(_05677_),
    .A3(_05686_),
    .Z(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12804_ (.A1(_05687_),
    .A2(_05688_),
    .ZN(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12805_ (.A1(_05675_),
    .A2(_05689_),
    .Z(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12806_ (.A1(_05657_),
    .A2(_05690_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12807_ (.I(_05610_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12808_ (.A1(_05606_),
    .A2(_05693_),
    .ZN(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12809_ (.A1(_05602_),
    .A2(_05611_),
    .B(_05694_),
    .ZN(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12810_ (.I(_05581_),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12811_ (.A1(_05696_),
    .A2(_05587_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12812_ (.A1(_05577_),
    .A2(_05578_),
    .B(_05588_),
    .ZN(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12813_ (.A1(_05697_),
    .A2(_05698_),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12814_ (.A1(_02762_),
    .A2(_00397_),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12815_ (.A1(_02854_),
    .A2(_00393_),
    .ZN(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12816_ (.A1(_02938_),
    .A2(_00390_),
    .ZN(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12817_ (.A1(_05701_),
    .A2(_05703_),
    .Z(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12818_ (.A1(_05700_),
    .A2(_05704_),
    .Z(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12819_ (.A1(_05608_),
    .A2(_05609_),
    .Z(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12820_ (.A1(_05608_),
    .A2(_05609_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12821_ (.A1(_05607_),
    .A2(_05706_),
    .B(_05707_),
    .ZN(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12822_ (.A1(_02940_),
    .A2(_00387_),
    .ZN(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12823_ (.A1(_03018_),
    .A2(_00384_),
    .ZN(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12824_ (.A1(_03189_),
    .A2(_00381_),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12825_ (.A1(_05709_),
    .A2(_05710_),
    .A3(_05711_),
    .Z(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12826_ (.A1(_05708_),
    .A2(_05712_),
    .Z(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12827_ (.A1(_05705_),
    .A2(_05714_),
    .Z(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12828_ (.A1(_05695_),
    .A2(_05699_),
    .A3(_05715_),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12829_ (.A1(_05692_),
    .A2(_05716_),
    .Z(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12830_ (.A1(_05654_),
    .A2(_05717_),
    .ZN(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12831_ (.A1(_05651_),
    .A2(_05718_),
    .ZN(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12832_ (.A1(_05641_),
    .A2(_05643_),
    .A3(_05719_),
    .Z(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12833_ (.A1(_05546_),
    .A2(_05617_),
    .ZN(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12834_ (.A1(_05544_),
    .A2(_05618_),
    .B(_05721_),
    .ZN(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12835_ (.A1(_05720_),
    .A2(_05722_),
    .ZN(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12836_ (.A1(_05619_),
    .A2(_05622_),
    .ZN(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12837_ (.A1(_05623_),
    .A2(_05630_),
    .B(_05725_),
    .ZN(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12838_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-10] ),
    .A2(_05723_),
    .A3(_05726_),
    .Z(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12839_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-11] ),
    .A2(_05631_),
    .ZN(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12840_ (.A1(_05728_),
    .A2(_05639_),
    .ZN(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12841_ (.A1(_05727_),
    .A2(_05729_),
    .Z(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12842_ (.A1(_05280_),
    .A2(net30),
    .ZN(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12843_ (.A1(_05822_),
    .A2(_05730_),
    .B(_05731_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12844_ (.A1(_05822_),
    .A2(net31),
    .ZN(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12845_ (.A1(_05632_),
    .A2(_05727_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _12846_ (.A1(_05447_),
    .A2(_05537_),
    .A3(_05733_),
    .Z(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12847_ (.A1(_05723_),
    .A2(_05726_),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12848_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-10] ),
    .A2(_05736_),
    .ZN(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12849_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-10] ),
    .A2(_05736_),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12850_ (.A1(_05728_),
    .A2(_05737_),
    .B(_05738_),
    .ZN(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _12851_ (.A1(_05636_),
    .A2(_05733_),
    .B1(_05735_),
    .B2(_05360_),
    .C(_05739_),
    .ZN(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12852_ (.A1(_05648_),
    .A2(_05649_),
    .B(_05646_),
    .ZN(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12853_ (.A1(_05654_),
    .A2(_05717_),
    .ZN(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12854_ (.A1(_05651_),
    .A2(_05718_),
    .B(_05742_),
    .ZN(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12855_ (.A1(_05699_),
    .A2(_05715_),
    .Z(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12856_ (.A1(_05699_),
    .A2(_05715_),
    .Z(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12857_ (.A1(_05695_),
    .A2(_05744_),
    .B(_05746_),
    .ZN(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12858_ (.A1(_05701_),
    .A2(_05703_),
    .Z(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12859_ (.A1(_02762_),
    .A2(_00397_),
    .A3(_05704_),
    .ZN(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12860_ (.A1(_05748_),
    .A2(_05749_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12861_ (.A1(_05747_),
    .A2(_05750_),
    .Z(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12862_ (.A1(_05657_),
    .A2(_05690_),
    .ZN(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12863_ (.A1(_05692_),
    .A2(_05716_),
    .B(_05752_),
    .ZN(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12864_ (.A1(_05662_),
    .A2(_05674_),
    .ZN(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12865_ (.A1(_05675_),
    .A2(_05689_),
    .ZN(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12866_ (.A1(_05754_),
    .A2(_05755_),
    .ZN(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12867_ (.A1(_05663_),
    .A2(_05667_),
    .Z(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12868_ (.A1(_05668_),
    .A2(_05673_),
    .B(_05758_),
    .ZN(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12869_ (.A1(net54),
    .A2(_03725_),
    .B1(_03727_),
    .B2(net66),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12870_ (.A1(net66),
    .A2(net54),
    .A3(_03725_),
    .A4(_03727_),
    .ZN(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12871_ (.A1(_05760_),
    .A2(_05666_),
    .B(_05761_),
    .ZN(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12872_ (.I(_05762_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12873_ (.A1(net66),
    .A2(net54),
    .B(_03727_),
    .ZN(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12874_ (.A1(net86),
    .A2(net54),
    .A3(_03727_),
    .Z(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12875_ (.A1(_05764_),
    .A2(_05765_),
    .ZN(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12876_ (.A1(net70),
    .A2(_03725_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12877_ (.A1(_05766_),
    .A2(_05768_),
    .Z(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12878_ (.A1(_05763_),
    .A2(_05769_),
    .Z(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12879_ (.A1(_03556_),
    .A2(_00369_),
    .ZN(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12880_ (.A1(_00365_),
    .A2(_03558_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12881_ (.A1(_00361_),
    .A2(_03679_),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12882_ (.A1(_05771_),
    .A2(_05772_),
    .A3(_05773_),
    .Z(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12883_ (.I(_05774_),
    .ZN(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12884_ (.A1(_05770_),
    .A2(_05775_),
    .Z(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12885_ (.A1(_05759_),
    .A2(_05776_),
    .Z(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12886_ (.A1(_05683_),
    .A2(_05684_),
    .Z(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12887_ (.A1(_05683_),
    .A2(_05684_),
    .Z(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12888_ (.A1(_05682_),
    .A2(_05779_),
    .B(_05780_),
    .ZN(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12889_ (.A1(_05671_),
    .A2(_05672_),
    .Z(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12890_ (.A1(_05671_),
    .A2(_05672_),
    .Z(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12891_ (.A1(_05670_),
    .A2(_05782_),
    .B(_05783_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12892_ (.A1(_03340_),
    .A2(_00378_),
    .ZN(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12893_ (.A1(net147),
    .A2(_00375_),
    .ZN(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12894_ (.A1(_03485_),
    .A2(_00372_),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12895_ (.A1(_05785_),
    .A2(_05786_),
    .A3(_05787_),
    .Z(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12896_ (.A1(_05784_),
    .A2(_05788_),
    .Z(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12897_ (.I(_05790_),
    .ZN(_05791_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12898_ (.A1(_05781_),
    .A2(_05791_),
    .Z(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12899_ (.A1(_05777_),
    .A2(_05792_),
    .Z(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12900_ (.A1(_05757_),
    .A2(_05793_),
    .ZN(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12901_ (.I(_05712_),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12902_ (.A1(_05708_),
    .A2(_05795_),
    .ZN(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12903_ (.A1(_05705_),
    .A2(_05714_),
    .B(_05796_),
    .ZN(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12904_ (.I(_05681_),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12905_ (.I(_05687_),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12906_ (.A1(_05798_),
    .A2(_05685_),
    .B(_05799_),
    .ZN(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12907_ (.A1(_02854_),
    .A2(_00397_),
    .ZN(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12908_ (.A1(_02938_),
    .A2(_00393_),
    .ZN(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12909_ (.A1(_02940_),
    .A2(_00390_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12910_ (.A1(_05803_),
    .A2(_05804_),
    .Z(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12911_ (.A1(_05802_),
    .A2(_05805_),
    .Z(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12912_ (.A1(_05710_),
    .A2(_05711_),
    .Z(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12913_ (.A1(_05710_),
    .A2(_05711_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12914_ (.A1(_05709_),
    .A2(_05807_),
    .B(_05808_),
    .ZN(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12915_ (.A1(_03018_),
    .A2(_00387_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12916_ (.A1(_03189_),
    .A2(_00384_),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12917_ (.A1(_03266_),
    .A2(_00381_),
    .ZN(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12918_ (.A1(_05810_),
    .A2(_05812_),
    .A3(_05813_),
    .Z(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12919_ (.A1(_05809_),
    .A2(_05814_),
    .Z(_05815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12920_ (.A1(_05806_),
    .A2(_05815_),
    .Z(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12921_ (.A1(_05797_),
    .A2(_05801_),
    .A3(_05816_),
    .ZN(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12922_ (.A1(_05794_),
    .A2(_05817_),
    .Z(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12923_ (.A1(_05753_),
    .A2(_05818_),
    .ZN(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12924_ (.A1(_05751_),
    .A2(_05819_),
    .ZN(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12925_ (.A1(_05743_),
    .A2(_05820_),
    .ZN(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12926_ (.A1(_05741_),
    .A2(_05821_),
    .Z(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12927_ (.I(_05719_),
    .ZN(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12928_ (.A1(_05643_),
    .A2(_05824_),
    .ZN(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12929_ (.A1(_05643_),
    .A2(_05719_),
    .ZN(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12930_ (.A1(_05641_),
    .A2(_05826_),
    .ZN(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12931_ (.A1(_05825_),
    .A2(_05827_),
    .ZN(_05828_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12932_ (.A1(_05823_),
    .A2(_05828_),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12933_ (.A1(_05270_),
    .A2(_05439_),
    .ZN(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12934_ (.A1(_05623_),
    .A2(_05723_),
    .ZN(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12935_ (.A1(_05626_),
    .A2(_05831_),
    .Z(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12936_ (.A1(_05830_),
    .A2(_05832_),
    .Z(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12937_ (.A1(_05443_),
    .A2(_05832_),
    .Z(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12938_ (.A1(_05720_),
    .A2(_05722_),
    .Z(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12939_ (.A1(_05629_),
    .A2(_05831_),
    .ZN(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12940_ (.A1(_05720_),
    .A2(_05722_),
    .Z(_05838_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _12941_ (.A1(_05725_),
    .A2(_05836_),
    .B(_05837_),
    .C(_05838_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _12942_ (.A1(_05336_),
    .A2(_05834_),
    .B(_05835_),
    .C(_05839_),
    .ZN(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12943_ (.A1(_05829_),
    .A2(_05840_),
    .Z(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12944_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-9] ),
    .A2(_05841_),
    .ZN(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12945_ (.A1(_05740_),
    .A2(_05842_),
    .ZN(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12946_ (.A1(_05740_),
    .A2(_05842_),
    .Z(_05845_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12947_ (.A1(_05387_),
    .A2(_05843_),
    .A3(_05845_),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12948_ (.A1(_05732_),
    .A2(_05846_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12949_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-9] ),
    .A2(_05841_),
    .ZN(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12950_ (.A1(_05847_),
    .A2(_05845_),
    .ZN(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12951_ (.I(_05820_),
    .ZN(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12952_ (.A1(_05743_),
    .A2(_05849_),
    .ZN(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12953_ (.A1(_05741_),
    .A2(_05821_),
    .ZN(_05851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12954_ (.A1(_05748_),
    .A2(_05749_),
    .B(_05747_),
    .ZN(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12955_ (.A1(_05753_),
    .A2(_05818_),
    .ZN(_05853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12956_ (.A1(_05751_),
    .A2(_05819_),
    .B(_05853_),
    .ZN(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12957_ (.A1(_05801_),
    .A2(_05816_),
    .Z(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12958_ (.A1(_05801_),
    .A2(_05816_),
    .Z(_05856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12959_ (.A1(_05797_),
    .A2(_05855_),
    .B(_05856_),
    .ZN(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12960_ (.A1(_05803_),
    .A2(_05804_),
    .Z(_05858_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12961_ (.A1(_02854_),
    .A2(_00397_),
    .A3(_05805_),
    .ZN(_05859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12962_ (.A1(_05858_),
    .A2(_05859_),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12963_ (.A1(_05857_),
    .A2(_05860_),
    .Z(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12964_ (.A1(_05757_),
    .A2(_05793_),
    .ZN(_05862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12965_ (.A1(_05794_),
    .A2(_05817_),
    .B(_05862_),
    .ZN(_05863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12966_ (.A1(_05759_),
    .A2(_05776_),
    .ZN(_05865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12967_ (.A1(_05777_),
    .A2(_05792_),
    .ZN(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12968_ (.A1(_05865_),
    .A2(_05866_),
    .ZN(_05867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12969_ (.A1(_05770_),
    .A2(_05775_),
    .ZN(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12970_ (.A1(_05763_),
    .A2(_05769_),
    .B(_05868_),
    .ZN(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12971_ (.A1(_00369_),
    .A2(_03558_),
    .ZN(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12972_ (.A1(_00365_),
    .A2(_03679_),
    .ZN(_05871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12973_ (.A1(_00361_),
    .A2(_03725_),
    .ZN(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12974_ (.A1(_05870_),
    .A2(_05871_),
    .A3(_05872_),
    .Z(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12975_ (.A1(net70),
    .A2(_03725_),
    .B(_05764_),
    .ZN(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _12976_ (.A1(_05765_),
    .A2(_05874_),
    .B(net70),
    .C(_03727_),
    .ZN(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12977_ (.A1(net70),
    .A2(_03727_),
    .ZN(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12978_ (.A1(_05764_),
    .A2(_05877_),
    .ZN(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12979_ (.A1(_05876_),
    .A2(_05878_),
    .ZN(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12980_ (.A1(_05873_),
    .A2(_05879_),
    .Z(_05880_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12981_ (.A1(_05869_),
    .A2(_05880_),
    .Z(_05881_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12982_ (.A1(_05786_),
    .A2(_05787_),
    .Z(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12983_ (.A1(_05786_),
    .A2(_05787_),
    .Z(_05883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12984_ (.A1(_05785_),
    .A2(_05882_),
    .B(_05883_),
    .ZN(_05884_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12985_ (.A1(_05772_),
    .A2(_05773_),
    .Z(_05885_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12986_ (.A1(_05772_),
    .A2(_05773_),
    .Z(_05887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12987_ (.A1(_05771_),
    .A2(_05885_),
    .B(_05887_),
    .ZN(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12988_ (.A1(net147),
    .A2(_00378_),
    .ZN(_05889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12989_ (.A1(_03485_),
    .A2(_00375_),
    .ZN(_05890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12990_ (.A1(_03556_),
    .A2(_00372_),
    .ZN(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12991_ (.A1(_05889_),
    .A2(_05890_),
    .A3(_05891_),
    .Z(_05892_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12992_ (.A1(_05888_),
    .A2(_05892_),
    .Z(_05893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12993_ (.I(_05893_),
    .ZN(_05894_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12994_ (.A1(_05884_),
    .A2(_05894_),
    .Z(_05895_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12995_ (.A1(_05881_),
    .A2(_05895_),
    .Z(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12996_ (.A1(_05867_),
    .A2(_05896_),
    .ZN(_05898_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12997_ (.I(_05814_),
    .ZN(_05899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12998_ (.A1(_05809_),
    .A2(_05899_),
    .ZN(_05900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12999_ (.A1(_05806_),
    .A2(_05815_),
    .B(_05900_),
    .ZN(_05901_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13000_ (.I(_05784_),
    .ZN(_05902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13001_ (.A1(_05781_),
    .A2(_05791_),
    .ZN(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13002_ (.A1(_05902_),
    .A2(_05788_),
    .B(_05903_),
    .ZN(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13003_ (.A1(_02938_),
    .A2(_00397_),
    .ZN(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13004_ (.A1(_02940_),
    .A2(_00393_),
    .ZN(_05906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13005_ (.A1(_03018_),
    .A2(_00390_),
    .ZN(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13006_ (.A1(_05906_),
    .A2(_05907_),
    .Z(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13007_ (.A1(_05905_),
    .A2(_05909_),
    .Z(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13008_ (.A1(_05812_),
    .A2(_05813_),
    .Z(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13009_ (.A1(_05812_),
    .A2(_05813_),
    .Z(_05912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13010_ (.A1(_05810_),
    .A2(_05911_),
    .B(_05912_),
    .ZN(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13011_ (.A1(_03189_),
    .A2(_00387_),
    .ZN(_05914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13012_ (.A1(_03266_),
    .A2(_00384_),
    .ZN(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13013_ (.A1(_03340_),
    .A2(_00381_),
    .ZN(_05916_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13014_ (.A1(_05914_),
    .A2(_05915_),
    .A3(_05916_),
    .Z(_05917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13015_ (.A1(_05913_),
    .A2(_05917_),
    .Z(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13016_ (.A1(_05910_),
    .A2(_05918_),
    .Z(_05920_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13017_ (.A1(_05901_),
    .A2(_05904_),
    .A3(_05920_),
    .ZN(_05921_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13018_ (.A1(_05898_),
    .A2(_05921_),
    .Z(_05922_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13019_ (.A1(_05863_),
    .A2(_05922_),
    .ZN(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13020_ (.A1(_05861_),
    .A2(_05923_),
    .ZN(_05924_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13021_ (.A1(_05852_),
    .A2(_05854_),
    .A3(_05924_),
    .Z(_05925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13022_ (.A1(_05850_),
    .A2(_05851_),
    .B(_05925_),
    .ZN(_05926_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13023_ (.A1(_05850_),
    .A2(_05851_),
    .A3(_05925_),
    .Z(_05927_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13024_ (.A1(_05926_),
    .A2(_05927_),
    .Z(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13025_ (.A1(_05823_),
    .A2(_05828_),
    .ZN(_05929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13026_ (.A1(_05829_),
    .A2(_05840_),
    .B(_05929_),
    .ZN(_05931_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13027_ (.A1(_05928_),
    .A2(_05931_),
    .ZN(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13028_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-8] ),
    .A2(_05932_),
    .ZN(_05933_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13029_ (.A1(_05848_),
    .A2(_05933_),
    .Z(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13030_ (.A1(_05280_),
    .A2(net32),
    .ZN(_05935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13031_ (.A1(_05822_),
    .A2(_05934_),
    .B(_05935_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13032_ (.A1(_05858_),
    .A2(_05859_),
    .B(_05857_),
    .ZN(_05936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13033_ (.A1(_05863_),
    .A2(_05922_),
    .ZN(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13034_ (.A1(_05861_),
    .A2(_05923_),
    .B(_05937_),
    .ZN(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13035_ (.A1(_05904_),
    .A2(_05920_),
    .Z(_05939_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13036_ (.A1(_05904_),
    .A2(_05920_),
    .Z(_05941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13037_ (.A1(_05901_),
    .A2(_05939_),
    .B(_05941_),
    .ZN(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13038_ (.A1(_05906_),
    .A2(_05907_),
    .Z(_05943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13039_ (.A1(_02938_),
    .A2(_00397_),
    .A3(_05909_),
    .ZN(_05944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13040_ (.A1(_05943_),
    .A2(_05944_),
    .ZN(_05945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13041_ (.A1(_05942_),
    .A2(_05945_),
    .Z(_05946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13042_ (.A1(_05867_),
    .A2(_05896_),
    .ZN(_05947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13043_ (.A1(_05898_),
    .A2(_05921_),
    .B(_05947_),
    .ZN(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13044_ (.A1(_05869_),
    .A2(_05880_),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13045_ (.A1(_05881_),
    .A2(_05895_),
    .ZN(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13046_ (.A1(_05949_),
    .A2(_05950_),
    .ZN(_05952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13047_ (.A1(net70),
    .A2(_05765_),
    .ZN(_05953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13048_ (.A1(_05873_),
    .A2(_05879_),
    .B(_05953_),
    .ZN(_05954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13049_ (.A1(_00369_),
    .A2(_03679_),
    .ZN(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13050_ (.A1(_00365_),
    .A2(_03725_),
    .ZN(_05956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13051_ (.A1(_00361_),
    .A2(_03727_),
    .ZN(_05957_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13052_ (.A1(_05955_),
    .A2(_05956_),
    .A3(_05957_),
    .Z(_05958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13053_ (.A1(_05878_),
    .A2(_05953_),
    .ZN(_05959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13054_ (.A1(_05958_),
    .A2(_05959_),
    .Z(_05960_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13055_ (.A1(_05954_),
    .A2(_05960_),
    .Z(_05961_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13056_ (.A1(_05890_),
    .A2(_05891_),
    .Z(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13057_ (.A1(_05890_),
    .A2(_05891_),
    .Z(_05964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13058_ (.A1(_05889_),
    .A2(_05963_),
    .B(_05964_),
    .ZN(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13059_ (.A1(_05871_),
    .A2(_05872_),
    .Z(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13060_ (.A1(_05871_),
    .A2(_05872_),
    .Z(_05967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13061_ (.A1(_05870_),
    .A2(_05966_),
    .B(_05967_),
    .ZN(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13062_ (.A1(_03485_),
    .A2(_00378_),
    .ZN(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13063_ (.A1(_03556_),
    .A2(_00375_),
    .ZN(_05970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13064_ (.A1(_00372_),
    .A2(_03558_),
    .ZN(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13065_ (.A1(_05969_),
    .A2(_05970_),
    .A3(_05971_),
    .Z(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13066_ (.A1(_05968_),
    .A2(_05972_),
    .Z(_05974_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13067_ (.I(_05974_),
    .ZN(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13068_ (.A1(_05965_),
    .A2(_05975_),
    .Z(_05976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13069_ (.A1(_05961_),
    .A2(_05976_),
    .Z(_05977_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13070_ (.A1(_05952_),
    .A2(_05977_),
    .ZN(_05978_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13071_ (.I(_05917_),
    .ZN(_05979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13072_ (.A1(_05913_),
    .A2(_05979_),
    .ZN(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13073_ (.A1(_05910_),
    .A2(_05918_),
    .B(_05980_),
    .ZN(_05981_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13074_ (.I(_05888_),
    .ZN(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13075_ (.A1(_05884_),
    .A2(_05894_),
    .ZN(_05983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13076_ (.A1(_05982_),
    .A2(_05892_),
    .B(_05983_),
    .ZN(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13077_ (.A1(_02940_),
    .A2(_00397_),
    .ZN(_05986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13078_ (.A1(_03018_),
    .A2(_00393_),
    .ZN(_05987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13079_ (.A1(_03189_),
    .A2(_00390_),
    .ZN(_05988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13080_ (.A1(_05987_),
    .A2(_05988_),
    .Z(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13081_ (.A1(_05986_),
    .A2(_05989_),
    .Z(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13082_ (.A1(_05915_),
    .A2(_05916_),
    .Z(_05991_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13083_ (.A1(_05915_),
    .A2(_05916_),
    .Z(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13084_ (.A1(_05914_),
    .A2(_05991_),
    .B(_05992_),
    .ZN(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13085_ (.A1(_03266_),
    .A2(_00387_),
    .ZN(_05994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13086_ (.A1(_03340_),
    .A2(_00384_),
    .ZN(_05996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13087_ (.A1(net147),
    .A2(_00381_),
    .ZN(_05997_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13088_ (.A1(_05994_),
    .A2(_05996_),
    .A3(_05997_),
    .Z(_05998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13089_ (.A1(_05993_),
    .A2(_05998_),
    .Z(_05999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13090_ (.A1(_05990_),
    .A2(_05999_),
    .Z(_06000_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13091_ (.A1(_05981_),
    .A2(_05985_),
    .A3(_06000_),
    .ZN(_06001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13092_ (.A1(_05978_),
    .A2(_06001_),
    .Z(_06002_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13093_ (.A1(_05948_),
    .A2(_06002_),
    .ZN(_06003_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13094_ (.A1(_05946_),
    .A2(_06003_),
    .ZN(_06004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13095_ (.I(_06004_),
    .ZN(_06005_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13096_ (.A1(_05938_),
    .A2(_06005_),
    .Z(_06007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13097_ (.A1(_05936_),
    .A2(_06007_),
    .Z(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13098_ (.I(_05924_),
    .ZN(_06009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13099_ (.A1(_05854_),
    .A2(_06009_),
    .ZN(_06010_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13100_ (.A1(_05854_),
    .A2(_06009_),
    .Z(_06011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13101_ (.A1(_05852_),
    .A2(_06010_),
    .A3(_06011_),
    .ZN(_06012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13102_ (.A1(_06010_),
    .A2(_06012_),
    .ZN(_06013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13103_ (.A1(_06008_),
    .A2(_06013_),
    .Z(_06014_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _13104_ (.I(_06014_),
    .ZN(_06015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13105_ (.A1(_05830_),
    .A2(_05832_),
    .ZN(_06016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13106_ (.A1(_05443_),
    .A2(_05832_),
    .ZN(_06018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13107_ (.A1(_05725_),
    .A2(_05836_),
    .B(_05838_),
    .ZN(_06019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13108_ (.A1(_05629_),
    .A2(_05831_),
    .B(_06019_),
    .ZN(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _13109_ (.A1(_05250_),
    .A2(_06016_),
    .B(_06018_),
    .C(_06020_),
    .ZN(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13110_ (.A1(_05829_),
    .A2(_05928_),
    .ZN(_06022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13111_ (.A1(_05823_),
    .A2(_05828_),
    .Z(_06023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13112_ (.A1(_06023_),
    .A2(_05926_),
    .ZN(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13113_ (.A1(_05927_),
    .A2(_06024_),
    .ZN(_06025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13114_ (.A1(_06021_),
    .A2(_06022_),
    .B(_06025_),
    .ZN(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13115_ (.A1(_06015_),
    .A2(_06026_),
    .Z(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13116_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-7] ),
    .A2(_06027_),
    .Z(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13117_ (.I(_06029_),
    .ZN(_06030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13118_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-8] ),
    .A2(_05932_),
    .ZN(_06031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13119_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-8] ),
    .A2(_05932_),
    .ZN(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13120_ (.A1(_05847_),
    .A2(_06031_),
    .B(_06032_),
    .ZN(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13121_ (.A1(_05842_),
    .A2(_05933_),
    .Z(_06034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13122_ (.A1(net77),
    .A2(_06034_),
    .ZN(_06035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13123_ (.A1(_06033_),
    .A2(_06035_),
    .ZN(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13124_ (.A1(_06030_),
    .A2(_06036_),
    .ZN(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _13125_ (.A1(_06029_),
    .A2(_06033_),
    .A3(_06035_),
    .B(_05182_),
    .ZN(_06038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13126_ (.A1(_05280_),
    .A2(net33),
    .ZN(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13127_ (.A1(_06037_),
    .A2(_06038_),
    .B(_06040_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13128_ (.A1(_05943_),
    .A2(_05944_),
    .B(_05942_),
    .ZN(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13129_ (.A1(_05948_),
    .A2(_06002_),
    .ZN(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13130_ (.A1(_05946_),
    .A2(_06003_),
    .B(_06042_),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13131_ (.A1(_05985_),
    .A2(_06000_),
    .Z(_06044_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13132_ (.A1(_05985_),
    .A2(_06000_),
    .Z(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13133_ (.A1(_05981_),
    .A2(_06044_),
    .B(_06045_),
    .ZN(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13134_ (.A1(_05987_),
    .A2(_05988_),
    .Z(_06047_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13135_ (.A1(_02940_),
    .A2(_00397_),
    .A3(_05989_),
    .ZN(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13136_ (.A1(_06047_),
    .A2(_06048_),
    .ZN(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13137_ (.A1(_06046_),
    .A2(_06049_),
    .Z(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13138_ (.A1(_05952_),
    .A2(_05977_),
    .ZN(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13139_ (.A1(_05978_),
    .A2(_06001_),
    .B(_06051_),
    .ZN(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13140_ (.A1(_05954_),
    .A2(_05960_),
    .ZN(_06053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13141_ (.A1(_05961_),
    .A2(_05976_),
    .ZN(_06054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13142_ (.A1(_06053_),
    .A2(_06054_),
    .ZN(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13143_ (.A1(_05958_),
    .A2(_05959_),
    .B(_05953_),
    .ZN(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13144_ (.A1(_00369_),
    .A2(_03725_),
    .ZN(_06057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13145_ (.A1(_00365_),
    .A2(_03727_),
    .ZN(_06058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13146_ (.A1(_05957_),
    .A2(_06058_),
    .Z(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13147_ (.A1(_06057_),
    .A2(_06060_),
    .Z(_06061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13148_ (.A1(_05959_),
    .A2(_06061_),
    .Z(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13149_ (.A1(_06056_),
    .A2(_06062_),
    .Z(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13150_ (.A1(_05970_),
    .A2(_05971_),
    .Z(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13151_ (.A1(_05970_),
    .A2(_05971_),
    .Z(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13152_ (.A1(_05969_),
    .A2(_06064_),
    .B(_06065_),
    .ZN(_06066_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13153_ (.A1(_05956_),
    .A2(_05957_),
    .Z(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13154_ (.A1(_05956_),
    .A2(_05957_),
    .Z(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13155_ (.A1(_05955_),
    .A2(_06067_),
    .B(_06068_),
    .ZN(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13156_ (.A1(_03556_),
    .A2(_00378_),
    .ZN(_06071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13157_ (.A1(_00375_),
    .A2(_03558_),
    .ZN(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13158_ (.A1(_00372_),
    .A2(_03679_),
    .ZN(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13159_ (.A1(_06071_),
    .A2(_06072_),
    .A3(_06073_),
    .Z(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13160_ (.A1(_06069_),
    .A2(_06074_),
    .Z(_06075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13161_ (.I(_06075_),
    .ZN(_06076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13162_ (.A1(_06066_),
    .A2(_06076_),
    .Z(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13163_ (.A1(_06063_),
    .A2(_06077_),
    .Z(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13164_ (.A1(_06055_),
    .A2(_06078_),
    .ZN(_06079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13165_ (.I(_05998_),
    .ZN(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13166_ (.A1(_05993_),
    .A2(_06080_),
    .ZN(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13167_ (.A1(_05990_),
    .A2(_05999_),
    .B(_06082_),
    .ZN(_06083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13168_ (.I(_05968_),
    .ZN(_06084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13169_ (.A1(_05965_),
    .A2(_05975_),
    .ZN(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13170_ (.A1(_06084_),
    .A2(_05972_),
    .B(_06085_),
    .ZN(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13171_ (.A1(_03018_),
    .A2(_00397_),
    .ZN(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13172_ (.A1(_03189_),
    .A2(_00393_),
    .ZN(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13173_ (.A1(_03266_),
    .A2(_00390_),
    .ZN(_06089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13174_ (.A1(_06088_),
    .A2(_06089_),
    .Z(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13175_ (.A1(_06087_),
    .A2(_06090_),
    .Z(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13176_ (.A1(_05996_),
    .A2(_05997_),
    .Z(_06093_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13177_ (.A1(_05996_),
    .A2(_05997_),
    .Z(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13178_ (.A1(_05994_),
    .A2(_06093_),
    .B(_06094_),
    .ZN(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13179_ (.A1(_03340_),
    .A2(_00387_),
    .ZN(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13180_ (.A1(net147),
    .A2(_00384_),
    .ZN(_06097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13181_ (.A1(_03485_),
    .A2(_00381_),
    .ZN(_06098_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13182_ (.A1(_06096_),
    .A2(_06097_),
    .A3(_06098_),
    .Z(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13183_ (.A1(_06095_),
    .A2(_06099_),
    .Z(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13184_ (.A1(_06091_),
    .A2(_06100_),
    .Z(_06101_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13185_ (.A1(_06083_),
    .A2(_06086_),
    .A3(_06101_),
    .ZN(_06102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13186_ (.A1(_06079_),
    .A2(_06102_),
    .Z(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13187_ (.A1(_06052_),
    .A2(_06104_),
    .ZN(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13188_ (.A1(_06050_),
    .A2(_06105_),
    .ZN(_06106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13189_ (.I(_06106_),
    .ZN(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13190_ (.A1(_06043_),
    .A2(_06107_),
    .Z(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13191_ (.A1(_06041_),
    .A2(_06108_),
    .ZN(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13192_ (.A1(_05938_),
    .A2(_06005_),
    .ZN(_06110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13193_ (.A1(_05936_),
    .A2(_06007_),
    .ZN(_06111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13194_ (.A1(_06110_),
    .A2(_06111_),
    .ZN(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13195_ (.A1(_06109_),
    .A2(_06112_),
    .Z(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _13196_ (.A1(_05829_),
    .A2(_05840_),
    .A3(_05928_),
    .B1(_06024_),
    .B2(_05927_),
    .ZN(_06115_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13197_ (.A1(_06008_),
    .A2(_06013_),
    .Z(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13198_ (.A1(_06014_),
    .A2(_06115_),
    .B(_06116_),
    .ZN(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13199_ (.A1(_06113_),
    .A2(_06117_),
    .Z(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _13200_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-6] ),
    .A2(_06118_),
    .Z(_06119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13201_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-6] ),
    .A2(_06118_),
    .ZN(_06120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13202_ (.A1(_06119_),
    .A2(_06120_),
    .ZN(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13203_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-7] ),
    .A2(_06027_),
    .Z(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13204_ (.A1(_06122_),
    .A2(_06037_),
    .ZN(_06123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13205_ (.A1(_06121_),
    .A2(_06123_),
    .Z(_06124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13206_ (.A1(_05280_),
    .A2(net34),
    .ZN(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13207_ (.A1(_05822_),
    .A2(_06124_),
    .B(_06126_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13208_ (.A1(_06029_),
    .A2(_06121_),
    .ZN(_06127_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13209_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-6] ),
    .A2(_06118_),
    .Z(_06128_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _13210_ (.A1(_06030_),
    .A2(_06119_),
    .A3(_06120_),
    .ZN(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _13211_ (.A1(_06122_),
    .A2(_06128_),
    .B1(_06129_),
    .B2(_06033_),
    .C(_06119_),
    .ZN(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _13212_ (.A1(_05740_),
    .A2(_06034_),
    .A3(_06127_),
    .B(_06130_),
    .ZN(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13213_ (.A1(_06047_),
    .A2(_06048_),
    .B(_06046_),
    .ZN(_06132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13214_ (.A1(_06052_),
    .A2(_06104_),
    .ZN(_06133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13215_ (.A1(_06050_),
    .A2(_06105_),
    .B(_06133_),
    .ZN(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13216_ (.A1(_06088_),
    .A2(_06089_),
    .Z(_06136_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13217_ (.A1(_03018_),
    .A2(_00397_),
    .A3(_06090_),
    .ZN(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13218_ (.A1(_06086_),
    .A2(_06101_),
    .Z(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13219_ (.A1(_06086_),
    .A2(_06101_),
    .Z(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13220_ (.A1(_06083_),
    .A2(_06138_),
    .B(_06139_),
    .ZN(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13221_ (.A1(_06136_),
    .A2(_06137_),
    .B(_06140_),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13222_ (.A1(_06136_),
    .A2(_06137_),
    .A3(_06140_),
    .Z(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13223_ (.A1(_06141_),
    .A2(_06142_),
    .ZN(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13224_ (.A1(_06055_),
    .A2(_06078_),
    .ZN(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13225_ (.A1(_06079_),
    .A2(_06102_),
    .B(_06144_),
    .ZN(_06145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13226_ (.A1(_06056_),
    .A2(_06062_),
    .ZN(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13227_ (.A1(_06063_),
    .A2(_06077_),
    .ZN(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13228_ (.A1(_06147_),
    .A2(_06148_),
    .ZN(_06149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13229_ (.A1(_05959_),
    .A2(_06061_),
    .B(_05953_),
    .ZN(_06150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13230_ (.A1(_00369_),
    .A2(_03727_),
    .ZN(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13231_ (.A1(_06060_),
    .A2(_06151_),
    .Z(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13232_ (.A1(_05959_),
    .A2(_06152_),
    .Z(_06153_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13233_ (.A1(_06150_),
    .A2(_06153_),
    .ZN(_06154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13234_ (.A1(_06072_),
    .A2(_06073_),
    .Z(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13235_ (.A1(_06072_),
    .A2(_06073_),
    .Z(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13236_ (.A1(_06071_),
    .A2(_06155_),
    .B(_06156_),
    .ZN(_06158_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13237_ (.A1(_00361_),
    .A2(_00365_),
    .A3(_03727_),
    .ZN(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13238_ (.A1(_00369_),
    .A2(_03725_),
    .A3(_06060_),
    .ZN(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13239_ (.A1(_06159_),
    .A2(_06160_),
    .Z(_06161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13240_ (.A1(_00378_),
    .A2(_03558_),
    .ZN(_06162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13241_ (.A1(_00375_),
    .A2(_03679_),
    .ZN(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13242_ (.A1(_00372_),
    .A2(_03725_),
    .ZN(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13243_ (.A1(_06163_),
    .A2(_06164_),
    .Z(_06165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13244_ (.A1(_06162_),
    .A2(_06165_),
    .Z(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13245_ (.A1(_06161_),
    .A2(_06166_),
    .ZN(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13246_ (.A1(_06158_),
    .A2(_06167_),
    .Z(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13247_ (.A1(_06154_),
    .A2(_06169_),
    .Z(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13248_ (.A1(_06149_),
    .A2(_06170_),
    .ZN(_06171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13249_ (.I(_06099_),
    .ZN(_06172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13250_ (.A1(_06095_),
    .A2(_06172_),
    .ZN(_06173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13251_ (.A1(_06091_),
    .A2(_06100_),
    .B(_06173_),
    .ZN(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13252_ (.I(_06069_),
    .ZN(_06175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13253_ (.A1(_06066_),
    .A2(_06076_),
    .ZN(_06176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13254_ (.A1(_06175_),
    .A2(_06074_),
    .B(_06176_),
    .ZN(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13255_ (.A1(_03189_),
    .A2(_00397_),
    .ZN(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13256_ (.A1(_03266_),
    .A2(_00393_),
    .ZN(_06180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13257_ (.A1(_03340_),
    .A2(_00390_),
    .ZN(_06181_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13258_ (.A1(_06180_),
    .A2(_06181_),
    .Z(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13259_ (.A1(_06178_),
    .A2(_06182_),
    .Z(_06183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13260_ (.A1(_06097_),
    .A2(_06098_),
    .Z(_06184_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13261_ (.A1(_06097_),
    .A2(_06098_),
    .Z(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13262_ (.A1(_06096_),
    .A2(_06184_),
    .B(_06185_),
    .ZN(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13263_ (.A1(net147),
    .A2(_00387_),
    .ZN(_06187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13264_ (.A1(_03485_),
    .A2(_00384_),
    .ZN(_06188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13265_ (.A1(_03556_),
    .A2(_00381_),
    .ZN(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13266_ (.A1(_06187_),
    .A2(_06188_),
    .A3(_06189_),
    .Z(_06191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13267_ (.A1(_06186_),
    .A2(_06191_),
    .Z(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13268_ (.A1(_06183_),
    .A2(_06192_),
    .Z(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13269_ (.A1(_06174_),
    .A2(_06177_),
    .A3(_06193_),
    .ZN(_06194_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13270_ (.A1(_06171_),
    .A2(_06194_),
    .Z(_06195_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13271_ (.A1(_06145_),
    .A2(_06195_),
    .ZN(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13272_ (.A1(_06143_),
    .A2(_06196_),
    .Z(_06197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13273_ (.I(_06197_),
    .ZN(_06198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13274_ (.A1(_06134_),
    .A2(_06198_),
    .Z(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13275_ (.A1(_06132_),
    .A2(_06199_),
    .Z(_06200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13276_ (.A1(_06043_),
    .A2(_06107_),
    .ZN(_06201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13277_ (.A1(_06041_),
    .A2(_06108_),
    .ZN(_06202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13278_ (.A1(_06201_),
    .A2(_06202_),
    .ZN(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13279_ (.A1(_06200_),
    .A2(_06203_),
    .Z(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13280_ (.A1(_06110_),
    .A2(_06111_),
    .B(_06109_),
    .ZN(_06205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13281_ (.A1(_06110_),
    .A2(_06111_),
    .A3(_06109_),
    .ZN(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13282_ (.A1(_06116_),
    .A2(_06205_),
    .B(_06206_),
    .ZN(_06207_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _13283_ (.A1(_06015_),
    .A2(_06026_),
    .A3(_06113_),
    .B(_06207_),
    .ZN(_06208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13284_ (.A1(_06204_),
    .A2(_06208_),
    .Z(_06209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13285_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-5] ),
    .A2(_06209_),
    .Z(_06210_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13286_ (.A1(_06131_),
    .A2(_06210_),
    .Z(_06212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13287_ (.A1(_06131_),
    .A2(_06210_),
    .B(_05182_),
    .ZN(_06213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13288_ (.A1(_05280_),
    .A2(net35),
    .ZN(_06214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13289_ (.A1(_06212_),
    .A2(_06213_),
    .B(_06214_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13290_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-5] ),
    .A2(_06209_),
    .Z(_06215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13291_ (.A1(_06215_),
    .A2(_06212_),
    .ZN(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13292_ (.A1(_06134_),
    .A2(_06198_),
    .ZN(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13293_ (.A1(_06132_),
    .A2(_06199_),
    .ZN(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13294_ (.I(_06143_),
    .ZN(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13295_ (.A1(_06145_),
    .A2(_06195_),
    .ZN(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13296_ (.A1(_06219_),
    .A2(_06196_),
    .B(_06220_),
    .ZN(_06222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13297_ (.I(_06222_),
    .ZN(_06223_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13298_ (.A1(_06180_),
    .A2(_06181_),
    .Z(_06224_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13299_ (.A1(_03189_),
    .A2(_00397_),
    .A3(_06182_),
    .ZN(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13300_ (.A1(_06177_),
    .A2(_06193_),
    .Z(_06226_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13301_ (.A1(_06177_),
    .A2(_06193_),
    .Z(_06227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13302_ (.A1(_06174_),
    .A2(_06226_),
    .B(_06227_),
    .ZN(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13303_ (.A1(_06224_),
    .A2(_06225_),
    .B(_06228_),
    .ZN(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13304_ (.A1(_06224_),
    .A2(_06225_),
    .A3(_06228_),
    .Z(_06230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13305_ (.A1(_06229_),
    .A2(_06230_),
    .ZN(_06231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13306_ (.A1(_06149_),
    .A2(_06170_),
    .ZN(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13307_ (.A1(_06171_),
    .A2(_06194_),
    .B(_06233_),
    .ZN(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13308_ (.A1(_06150_),
    .A2(_06153_),
    .ZN(_06235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13309_ (.A1(_06154_),
    .A2(_06169_),
    .B(_06235_),
    .ZN(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _13310_ (.A1(_05953_),
    .A2(_06152_),
    .Z(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13311_ (.A1(_05953_),
    .A2(_05959_),
    .A3(_06152_),
    .ZN(_06238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _13312_ (.A1(_06237_),
    .A2(_06238_),
    .ZN(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13313_ (.A1(_00378_),
    .A2(_03558_),
    .A3(_06165_),
    .ZN(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13314_ (.A1(_06163_),
    .A2(_06164_),
    .B(_06240_),
    .ZN(_06241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13315_ (.A1(_00369_),
    .A2(_03727_),
    .A3(_06060_),
    .ZN(_06242_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _13316_ (.A1(_06159_),
    .A2(_06242_),
    .Z(_06244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13317_ (.A1(_00375_),
    .A2(_03725_),
    .ZN(_06245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13318_ (.A1(_00372_),
    .A2(_03727_),
    .ZN(_06246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13319_ (.A1(_06245_),
    .A2(_06246_),
    .ZN(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13320_ (.A1(_06245_),
    .A2(_06246_),
    .Z(_06248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13321_ (.A1(_06247_),
    .A2(_06248_),
    .ZN(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13322_ (.A1(_00378_),
    .A2(_03679_),
    .ZN(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13323_ (.A1(_06249_),
    .A2(_06250_),
    .ZN(_06251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13324_ (.A1(_06244_),
    .A2(_06251_),
    .Z(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13325_ (.A1(_06241_),
    .A2(_06252_),
    .ZN(_06253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13326_ (.A1(_06239_),
    .A2(_06253_),
    .Z(_06255_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13327_ (.A1(_06236_),
    .A2(_06255_),
    .ZN(_06256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13328_ (.I(_06191_),
    .ZN(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13329_ (.A1(_06186_),
    .A2(_06257_),
    .ZN(_06258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13330_ (.A1(_06183_),
    .A2(_06192_),
    .B(_06258_),
    .ZN(_06259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13331_ (.I(_06167_),
    .ZN(_06260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13332_ (.A1(_06158_),
    .A2(_06260_),
    .ZN(_06261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13333_ (.A1(_06161_),
    .A2(_06166_),
    .B(_06261_),
    .ZN(_06262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13334_ (.A1(_03266_),
    .A2(_00397_),
    .ZN(_06263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13335_ (.A1(_03340_),
    .A2(_00393_),
    .ZN(_06264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13336_ (.A1(net147),
    .A2(_00390_),
    .ZN(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13337_ (.A1(_06264_),
    .A2(_06266_),
    .Z(_06267_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13338_ (.A1(_06263_),
    .A2(_06267_),
    .Z(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13339_ (.I(_06268_),
    .ZN(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13340_ (.A1(_06188_),
    .A2(_06189_),
    .Z(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13341_ (.A1(_06188_),
    .A2(_06189_),
    .Z(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13342_ (.A1(_06187_),
    .A2(_06270_),
    .B(_06271_),
    .ZN(_06272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13343_ (.I(_06272_),
    .ZN(_06273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13344_ (.A1(_03485_),
    .A2(_00387_),
    .ZN(_06274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13345_ (.A1(_03556_),
    .A2(_00384_),
    .ZN(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13346_ (.A1(_00381_),
    .A2(_03558_),
    .ZN(_06277_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13347_ (.A1(_06274_),
    .A2(_06275_),
    .A3(_06277_),
    .Z(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13348_ (.A1(_06273_),
    .A2(_06278_),
    .Z(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13349_ (.A1(_06269_),
    .A2(_06279_),
    .Z(_06280_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13350_ (.A1(_06259_),
    .A2(_06262_),
    .A3(_06280_),
    .ZN(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13351_ (.A1(_06256_),
    .A2(_06281_),
    .Z(_06282_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13352_ (.A1(_06234_),
    .A2(_06282_),
    .ZN(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13353_ (.A1(_06231_),
    .A2(_06283_),
    .Z(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13354_ (.A1(_06223_),
    .A2(_06284_),
    .Z(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13355_ (.A1(_06141_),
    .A2(_06285_),
    .ZN(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13356_ (.A1(_06217_),
    .A2(_06218_),
    .B(_06286_),
    .ZN(_06288_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13357_ (.A1(_06217_),
    .A2(_06218_),
    .A3(_06286_),
    .Z(_06289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13358_ (.A1(_06288_),
    .A2(_06289_),
    .ZN(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13359_ (.A1(_06200_),
    .A2(_06203_),
    .Z(_06291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13360_ (.A1(_06204_),
    .A2(_06208_),
    .B(_06291_),
    .ZN(_06292_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13361_ (.A1(_06290_),
    .A2(_06292_),
    .ZN(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13362_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-4] ),
    .A2(_06293_),
    .Z(_06294_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13363_ (.A1(_06216_),
    .A2(_06294_),
    .Z(_06295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13364_ (.A1(_05280_),
    .A2(net21),
    .ZN(_06296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13365_ (.A1(_05822_),
    .A2(_06295_),
    .B(_06296_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13366_ (.A1(_05822_),
    .A2(net22),
    .ZN(_06298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13367_ (.I(_06289_),
    .ZN(_06299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13368_ (.A1(_06291_),
    .A2(_06288_),
    .B(_06299_),
    .ZN(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13369_ (.A1(_06204_),
    .A2(_06208_),
    .A3(_06290_),
    .ZN(_06301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13370_ (.A1(_06300_),
    .A2(_06301_),
    .ZN(_06302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13371_ (.A1(_06141_),
    .A2(_06285_),
    .ZN(_06303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13372_ (.A1(_06223_),
    .A2(_06284_),
    .B(_06303_),
    .ZN(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13373_ (.I(_06231_),
    .ZN(_06305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13374_ (.A1(_06234_),
    .A2(_06282_),
    .ZN(_06306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13375_ (.A1(_06305_),
    .A2(_06283_),
    .B(_06306_),
    .ZN(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13376_ (.A1(_06264_),
    .A2(_06266_),
    .Z(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13377_ (.A1(_03266_),
    .A2(_00397_),
    .A3(_06267_),
    .ZN(_06310_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13378_ (.A1(_06262_),
    .A2(_06280_),
    .Z(_06311_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13379_ (.A1(_06262_),
    .A2(_06280_),
    .Z(_06312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13380_ (.A1(_06259_),
    .A2(_06311_),
    .B(_06312_),
    .ZN(_06313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13381_ (.A1(_06309_),
    .A2(_06310_),
    .B(_06313_),
    .ZN(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13382_ (.A1(_06309_),
    .A2(_06310_),
    .A3(_06313_),
    .Z(_06315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13383_ (.A1(_06314_),
    .A2(_06315_),
    .ZN(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13384_ (.A1(_06236_),
    .A2(_06255_),
    .ZN(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13385_ (.A1(_06256_),
    .A2(_06281_),
    .B(_06317_),
    .ZN(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13386_ (.A1(_06239_),
    .A2(_06253_),
    .B(_06237_),
    .ZN(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13387_ (.A1(_06249_),
    .A2(_06250_),
    .B(_06248_),
    .ZN(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13388_ (.A1(_00372_),
    .A2(_00375_),
    .B(_03727_),
    .ZN(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13389_ (.A1(_00372_),
    .A2(_00375_),
    .A3(_03727_),
    .Z(_06323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13390_ (.A1(_06322_),
    .A2(_06323_),
    .ZN(_06324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13391_ (.A1(_00378_),
    .A2(_03725_),
    .ZN(_06325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13392_ (.A1(_06324_),
    .A2(_06325_),
    .Z(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13393_ (.A1(_06244_),
    .A2(_06326_),
    .Z(_06327_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13394_ (.A1(_06321_),
    .A2(_06327_),
    .ZN(_06328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13395_ (.A1(_06239_),
    .A2(_06328_),
    .Z(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13396_ (.A1(_06320_),
    .A2(_06329_),
    .Z(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13397_ (.I(_06330_),
    .ZN(_06331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13398_ (.A1(_06269_),
    .A2(_06279_),
    .ZN(_06332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13399_ (.A1(_06273_),
    .A2(_06278_),
    .B(_06332_),
    .ZN(_06333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13400_ (.A1(_06241_),
    .A2(_06252_),
    .ZN(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13401_ (.A1(_06244_),
    .A2(_06251_),
    .B(_06334_),
    .ZN(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13402_ (.A1(_03340_),
    .A2(_00397_),
    .ZN(_06336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13403_ (.A1(net147),
    .A2(_00393_),
    .ZN(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13404_ (.A1(_03485_),
    .A2(_00390_),
    .ZN(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13405_ (.A1(_06337_),
    .A2(_06338_),
    .Z(_06339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13406_ (.A1(_06336_),
    .A2(_06339_),
    .Z(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13407_ (.I(_06341_),
    .ZN(_06342_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13408_ (.A1(_06275_),
    .A2(_06277_),
    .Z(_06343_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13409_ (.A1(_06275_),
    .A2(_06277_),
    .Z(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13410_ (.A1(_06274_),
    .A2(_06343_),
    .B(_06344_),
    .ZN(_06345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13411_ (.I(_06345_),
    .ZN(_06346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13412_ (.A1(_03556_),
    .A2(_00387_),
    .ZN(_06347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13413_ (.A1(_00384_),
    .A2(_03558_),
    .ZN(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13414_ (.A1(_00381_),
    .A2(_03679_),
    .ZN(_06349_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13415_ (.A1(_06347_),
    .A2(_06348_),
    .A3(_06349_),
    .Z(_06350_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13416_ (.A1(_06346_),
    .A2(_06350_),
    .Z(_06352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13417_ (.A1(_06342_),
    .A2(_06352_),
    .Z(_06353_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13418_ (.A1(_06335_),
    .A2(_06353_),
    .Z(_06354_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13419_ (.A1(_06333_),
    .A2(_06354_),
    .ZN(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13420_ (.A1(_06331_),
    .A2(_06355_),
    .Z(_06356_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13421_ (.A1(_06318_),
    .A2(_06356_),
    .ZN(_06357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13422_ (.A1(_06316_),
    .A2(_06357_),
    .Z(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13423_ (.I(_06358_),
    .ZN(_06359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13424_ (.A1(_06307_),
    .A2(_06359_),
    .Z(_06360_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13425_ (.A1(_06229_),
    .A2(_06360_),
    .Z(_06361_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13426_ (.A1(_06304_),
    .A2(_06361_),
    .Z(_06363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13427_ (.A1(_06302_),
    .A2(_06363_),
    .Z(_06364_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13428_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-3] ),
    .A2(_06364_),
    .ZN(_06365_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13429_ (.A1(_06210_),
    .A2(_06294_),
    .Z(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13430_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-4] ),
    .A2(_06293_),
    .ZN(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13431_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-4] ),
    .A2(_06293_),
    .B(_06215_),
    .ZN(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13432_ (.A1(_06367_),
    .A2(_06368_),
    .ZN(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13433_ (.A1(_06131_),
    .A2(_06366_),
    .B(_06369_),
    .ZN(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13434_ (.A1(_06365_),
    .A2(_06370_),
    .ZN(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13435_ (.A1(_06365_),
    .A2(_06370_),
    .Z(_06372_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13436_ (.A1(_05387_),
    .A2(_06371_),
    .A3(_06372_),
    .ZN(_06374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13437_ (.A1(_06298_),
    .A2(_06374_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13438_ (.A1(_06304_),
    .A2(_06361_),
    .Z(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13439_ (.I(_06363_),
    .ZN(_06376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13440_ (.A1(_06300_),
    .A2(_06301_),
    .B(_06376_),
    .ZN(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13441_ (.A1(_06375_),
    .A2(_06377_),
    .ZN(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13442_ (.A1(_06307_),
    .A2(_06359_),
    .ZN(_06379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13443_ (.A1(_06229_),
    .A2(_06360_),
    .ZN(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13444_ (.A1(_06379_),
    .A2(_06380_),
    .ZN(_06381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13445_ (.I(_06316_),
    .ZN(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13446_ (.A1(_06318_),
    .A2(_06356_),
    .ZN(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13447_ (.A1(_06382_),
    .A2(_06357_),
    .B(_06384_),
    .ZN(_06385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13448_ (.A1(_06335_),
    .A2(_06353_),
    .ZN(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13449_ (.A1(_06333_),
    .A2(_06354_),
    .ZN(_06387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13450_ (.A1(_06386_),
    .A2(_06387_),
    .ZN(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13451_ (.A1(_03340_),
    .A2(_00397_),
    .A3(_06339_),
    .ZN(_06389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13452_ (.A1(_06337_),
    .A2(_06338_),
    .B(_06389_),
    .ZN(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13453_ (.A1(_06388_),
    .A2(_06390_),
    .Z(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13454_ (.A1(_06320_),
    .A2(_06329_),
    .ZN(_06392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13455_ (.A1(_06331_),
    .A2(_06355_),
    .B(_06392_),
    .ZN(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13456_ (.A1(_06239_),
    .A2(_06328_),
    .B(_06237_),
    .ZN(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _13457_ (.A1(_06322_),
    .A2(_06323_),
    .A3(_06325_),
    .ZN(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13458_ (.A1(_00378_),
    .A2(_03727_),
    .A3(_06324_),
    .ZN(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13459_ (.I(_06397_),
    .ZN(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13460_ (.A1(_00378_),
    .A2(_03727_),
    .B(_06324_),
    .ZN(_06399_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13461_ (.A1(_06398_),
    .A2(_06399_),
    .Z(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13462_ (.A1(_06244_),
    .A2(_06400_),
    .Z(_06401_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _13463_ (.A1(_06323_),
    .A2(_06396_),
    .A3(_06401_),
    .Z(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13464_ (.A1(_06323_),
    .A2(_06396_),
    .B(_06401_),
    .ZN(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13465_ (.A1(_06402_),
    .A2(_06403_),
    .ZN(_06404_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13466_ (.A1(_06239_),
    .A2(_06404_),
    .Z(_06406_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13467_ (.A1(_06395_),
    .A2(_06406_),
    .ZN(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13468_ (.A1(_06342_),
    .A2(_06352_),
    .ZN(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13469_ (.A1(_06346_),
    .A2(_06350_),
    .B(_06408_),
    .ZN(_06409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13470_ (.A1(_06321_),
    .A2(_06327_),
    .ZN(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13471_ (.A1(_06244_),
    .A2(_06326_),
    .B(_06410_),
    .ZN(_06411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13472_ (.A1(net147),
    .A2(_00397_),
    .ZN(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13473_ (.A1(_03485_),
    .A2(_00393_),
    .ZN(_06413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13474_ (.A1(_03556_),
    .A2(_00390_),
    .ZN(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13475_ (.A1(_06413_),
    .A2(_06414_),
    .Z(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13476_ (.A1(_06412_),
    .A2(_06415_),
    .Z(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13477_ (.I(_06417_),
    .ZN(_06418_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13478_ (.A1(_06348_),
    .A2(_06349_),
    .Z(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13479_ (.A1(_06348_),
    .A2(_06349_),
    .Z(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13480_ (.A1(_06347_),
    .A2(_06419_),
    .B(_06420_),
    .ZN(_06421_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13481_ (.I(_06421_),
    .ZN(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13482_ (.A1(_00387_),
    .A2(_03558_),
    .ZN(_06423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13483_ (.A1(_00384_),
    .A2(_03679_),
    .ZN(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13484_ (.A1(_00381_),
    .A2(_03725_),
    .ZN(_06425_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13485_ (.A1(_06423_),
    .A2(_06424_),
    .A3(_06425_),
    .Z(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13486_ (.A1(_06422_),
    .A2(_06426_),
    .Z(_06428_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13487_ (.A1(_06418_),
    .A2(_06428_),
    .Z(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13488_ (.A1(_06411_),
    .A2(_06429_),
    .Z(_06430_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13489_ (.A1(_06409_),
    .A2(_06430_),
    .ZN(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13490_ (.A1(_06407_),
    .A2(_06431_),
    .Z(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13491_ (.A1(_06393_),
    .A2(_06432_),
    .Z(_06433_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13492_ (.A1(_06391_),
    .A2(_06433_),
    .Z(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13493_ (.A1(_06385_),
    .A2(_06434_),
    .Z(_06435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13494_ (.A1(_06314_),
    .A2(_06435_),
    .Z(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13495_ (.A1(_06381_),
    .A2(_06436_),
    .Z(_06437_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13496_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ),
    .A2(_06378_),
    .A3(_06437_),
    .Z(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13497_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-3] ),
    .A2(_06364_),
    .ZN(_06439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13498_ (.A1(_06439_),
    .A2(_06372_),
    .ZN(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13499_ (.A1(_06438_),
    .A2(_06440_),
    .Z(_06441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13500_ (.A1(_05280_),
    .A2(net23),
    .ZN(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13501_ (.A1(_05822_),
    .A2(_06441_),
    .B(_06442_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13502_ (.A1(_06365_),
    .A2(_06438_),
    .ZN(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13503_ (.A1(_06210_),
    .A2(_06294_),
    .ZN(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _13504_ (.A1(_06365_),
    .A2(_06444_),
    .A3(_06438_),
    .ZN(_06445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13505_ (.A1(_06375_),
    .A2(_06377_),
    .B(_06437_),
    .ZN(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _13506_ (.A1(_06375_),
    .A2(_06377_),
    .A3(_06437_),
    .Z(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13507_ (.A1(_06446_),
    .A2(_06448_),
    .B(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ),
    .ZN(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13508_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ),
    .A2(_06446_),
    .A3(_06448_),
    .ZN(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13509_ (.A1(_06439_),
    .A2(_06449_),
    .B(_06450_),
    .ZN(_06451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _13510_ (.A1(_06369_),
    .A2(_06443_),
    .B1(_06445_),
    .B2(_06131_),
    .C(_06451_),
    .ZN(_06452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13511_ (.A1(_06381_),
    .A2(_06436_),
    .ZN(_06453_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13512_ (.A1(_06453_),
    .A2(_06446_),
    .Z(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13513_ (.A1(_06385_),
    .A2(_06434_),
    .ZN(_06455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13514_ (.A1(_06314_),
    .A2(_06435_),
    .ZN(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13515_ (.A1(_06455_),
    .A2(_06456_),
    .ZN(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13516_ (.A1(_06388_),
    .A2(_06390_),
    .Z(_06459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13517_ (.A1(_06393_),
    .A2(_06432_),
    .ZN(_06460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13518_ (.A1(_06391_),
    .A2(_06433_),
    .ZN(_06461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13519_ (.A1(_06460_),
    .A2(_06461_),
    .ZN(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13520_ (.A1(_06413_),
    .A2(_06414_),
    .Z(_06463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13521_ (.A1(net147),
    .A2(_00397_),
    .A3(_06415_),
    .ZN(_06464_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13522_ (.A1(_06411_),
    .A2(_06429_),
    .Z(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13523_ (.A1(_06409_),
    .A2(_06430_),
    .B(_06465_),
    .ZN(_06466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13524_ (.A1(_06463_),
    .A2(_06464_),
    .B(_06466_),
    .ZN(_06467_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13525_ (.A1(_06463_),
    .A2(_06464_),
    .A3(_06466_),
    .Z(_06468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13526_ (.A1(_06467_),
    .A2(_06468_),
    .ZN(_06470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13527_ (.A1(_06395_),
    .A2(_06406_),
    .ZN(_06471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13528_ (.A1(_06407_),
    .A2(_06431_),
    .B(_06471_),
    .ZN(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13529_ (.A1(_06239_),
    .A2(_06404_),
    .B(_06237_),
    .ZN(_06473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13530_ (.A1(_06323_),
    .A2(_06398_),
    .B(_06401_),
    .ZN(_06474_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _13531_ (.A1(_06323_),
    .A2(_06398_),
    .A3(_06401_),
    .Z(_06475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13532_ (.A1(_06474_),
    .A2(_06475_),
    .ZN(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13533_ (.A1(_06239_),
    .A2(_06476_),
    .Z(_06477_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13534_ (.A1(_06473_),
    .A2(_06477_),
    .ZN(_06478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13535_ (.A1(_06418_),
    .A2(_06428_),
    .ZN(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13536_ (.A1(_06422_),
    .A2(_06426_),
    .B(_06479_),
    .ZN(_06481_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13537_ (.A1(_06244_),
    .A2(_06400_),
    .Z(_06482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13538_ (.A1(_06482_),
    .A2(_06403_),
    .ZN(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13539_ (.A1(_03485_),
    .A2(_00397_),
    .ZN(_06484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13540_ (.A1(_03556_),
    .A2(_00393_),
    .ZN(_06485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13541_ (.A1(_00390_),
    .A2(_03558_),
    .ZN(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13542_ (.A1(_06485_),
    .A2(_06486_),
    .Z(_06487_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13543_ (.A1(_06484_),
    .A2(_06487_),
    .Z(_06488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13544_ (.A1(_06424_),
    .A2(_06425_),
    .Z(_06489_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13545_ (.A1(_06424_),
    .A2(_06425_),
    .Z(_06490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13546_ (.A1(_06423_),
    .A2(_06489_),
    .B(_06490_),
    .ZN(_06492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13547_ (.A1(_00384_),
    .A2(_03725_),
    .ZN(_06493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13548_ (.A1(_00381_),
    .A2(_03727_),
    .ZN(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13549_ (.A1(_00387_),
    .A2(_03679_),
    .ZN(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13550_ (.A1(_06493_),
    .A2(_06494_),
    .A3(_06495_),
    .Z(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13551_ (.A1(_06492_),
    .A2(_06496_),
    .Z(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13552_ (.A1(_06488_),
    .A2(_06497_),
    .Z(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13553_ (.A1(_06483_),
    .A2(_06498_),
    .Z(_06499_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13554_ (.A1(_06481_),
    .A2(_06499_),
    .ZN(_06500_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13555_ (.A1(_06478_),
    .A2(_06500_),
    .Z(_06501_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13556_ (.A1(_06472_),
    .A2(_06501_),
    .Z(_06503_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13557_ (.A1(_06470_),
    .A2(_06503_),
    .Z(_06504_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13558_ (.A1(_06462_),
    .A2(_06504_),
    .Z(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13559_ (.A1(_06459_),
    .A2(_06505_),
    .Z(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13560_ (.A1(_06457_),
    .A2(_06506_),
    .ZN(_06507_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13561_ (.A1(_06454_),
    .A2(_06507_),
    .Z(_06508_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13562_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-1] ),
    .A2(_06508_),
    .ZN(_06509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13563_ (.A1(_06452_),
    .A2(_06509_),
    .ZN(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _13564_ (.A1(_06452_),
    .A2(_06509_),
    .Z(_06511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13565_ (.A1(_06510_),
    .A2(_06511_),
    .ZN(_06512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13566_ (.A1(_05280_),
    .A2(net24),
    .ZN(_06514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13567_ (.A1(_05822_),
    .A2(_06512_),
    .B(_06514_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13568_ (.A1(_06457_),
    .A2(_06506_),
    .ZN(_06515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13569_ (.A1(_06454_),
    .A2(_06507_),
    .B(_06515_),
    .ZN(_06516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13570_ (.A1(_06462_),
    .A2(_06504_),
    .ZN(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13571_ (.A1(_06459_),
    .A2(_06505_),
    .ZN(_06518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13572_ (.A1(_06517_),
    .A2(_06518_),
    .ZN(_06519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13573_ (.A1(_06472_),
    .A2(_06501_),
    .ZN(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13574_ (.A1(_06470_),
    .A2(_06503_),
    .ZN(_06521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13575_ (.A1(_06520_),
    .A2(_06521_),
    .ZN(_06522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13576_ (.I(_06522_),
    .ZN(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13577_ (.A1(_06473_),
    .A2(_06477_),
    .ZN(_06525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13578_ (.A1(_06478_),
    .A2(_06500_),
    .B(_06525_),
    .ZN(_06526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13579_ (.A1(_06237_),
    .A2(_06476_),
    .ZN(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13580_ (.A1(_06237_),
    .A2(_06239_),
    .A3(_06476_),
    .Z(_06528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13581_ (.A1(_06527_),
    .A2(_06528_),
    .ZN(_06529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13582_ (.I(_06496_),
    .ZN(_06530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13583_ (.A1(_06492_),
    .A2(_06530_),
    .ZN(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13584_ (.A1(_06488_),
    .A2(_06497_),
    .B(_06531_),
    .ZN(_06532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13585_ (.A1(_06482_),
    .A2(_06474_),
    .ZN(_06533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13586_ (.A1(_03556_),
    .A2(_00397_),
    .ZN(_06535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13587_ (.A1(_00393_),
    .A2(_03558_),
    .ZN(_06536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13588_ (.A1(_00390_),
    .A2(_03679_),
    .ZN(_06537_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13589_ (.A1(_06535_),
    .A2(_06536_),
    .A3(_06537_),
    .Z(_06538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13590_ (.I(_06538_),
    .ZN(_06539_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13591_ (.A1(_06493_),
    .A2(_06494_),
    .Z(_06540_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13592_ (.A1(_06493_),
    .A2(_06494_),
    .Z(_06541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13593_ (.A1(_06540_),
    .A2(_06495_),
    .B(_06541_),
    .ZN(_06542_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13594_ (.I(_06542_),
    .ZN(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13595_ (.A1(_00387_),
    .A2(_03725_),
    .ZN(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13596_ (.A1(_00381_),
    .A2(_00384_),
    .B(_03727_),
    .ZN(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13597_ (.A1(_00381_),
    .A2(_00384_),
    .A3(_03727_),
    .Z(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13598_ (.A1(_06545_),
    .A2(_06546_),
    .ZN(_06547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13599_ (.A1(_06544_),
    .A2(_06547_),
    .Z(_06548_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13600_ (.A1(_06543_),
    .A2(_06548_),
    .Z(_06549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13601_ (.A1(_06539_),
    .A2(_06549_),
    .Z(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13602_ (.A1(_06532_),
    .A2(_06533_),
    .A3(_06550_),
    .ZN(_06551_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13603_ (.A1(_06529_),
    .A2(_06551_),
    .ZN(_06552_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13604_ (.A1(_06526_),
    .A2(_06552_),
    .ZN(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13605_ (.A1(_06483_),
    .A2(_06498_),
    .Z(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13606_ (.A1(_06481_),
    .A2(_06499_),
    .B(_06554_),
    .ZN(_06556_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13607_ (.A1(_06485_),
    .A2(_06486_),
    .Z(_06557_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13608_ (.A1(_03485_),
    .A2(_00397_),
    .A3(_06487_),
    .ZN(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13609_ (.A1(_06557_),
    .A2(_06558_),
    .ZN(_06559_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13610_ (.A1(_06556_),
    .A2(_06559_),
    .ZN(_06560_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13611_ (.A1(_06553_),
    .A2(_06560_),
    .Z(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13612_ (.A1(_06524_),
    .A2(_06561_),
    .Z(_06562_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13613_ (.A1(_06467_),
    .A2(_06562_),
    .Z(_06563_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13614_ (.A1(_06519_),
    .A2(_06563_),
    .Z(_06564_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13615_ (.A1(_06516_),
    .A2(_06564_),
    .Z(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13616_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-1] ),
    .A2(_06508_),
    .Z(_06567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13617_ (.I(_06567_),
    .ZN(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13618_ (.A1(_06568_),
    .A2(_06511_),
    .ZN(_06569_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13619_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[0] ),
    .A2(_06565_),
    .A3(_06569_),
    .Z(_06570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13620_ (.I0(net25),
    .I1(_06570_),
    .S(_05171_),
    .Z(_06571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13621_ (.I(_06571_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13622_ (.A1(_06519_),
    .A2(_06563_),
    .Z(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13623_ (.A1(_06516_),
    .A2(_06564_),
    .B(_06572_),
    .ZN(_06573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13624_ (.A1(_06467_),
    .A2(_06562_),
    .ZN(_06574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13625_ (.A1(_06524_),
    .A2(_06561_),
    .B(_06574_),
    .ZN(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13626_ (.I(_06528_),
    .ZN(_06577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13627_ (.A1(_06577_),
    .A2(_06551_),
    .B(_06527_),
    .ZN(_06578_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13628_ (.A1(_06533_),
    .A2(_06578_),
    .Z(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13629_ (.A1(_00387_),
    .A2(_03725_),
    .B(_06545_),
    .ZN(_06580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13630_ (.A1(_06546_),
    .A2(_06580_),
    .ZN(_06581_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13631_ (.I(_06560_),
    .ZN(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13632_ (.A1(_06526_),
    .A2(_06552_),
    .ZN(_06583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13633_ (.A1(_06553_),
    .A2(_06582_),
    .B(_06583_),
    .ZN(_06584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13634_ (.A1(_06557_),
    .A2(_06558_),
    .B(_06556_),
    .ZN(_06585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13635_ (.A1(_00393_),
    .A2(_03679_),
    .ZN(_06586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13636_ (.A1(_00390_),
    .A2(_03725_),
    .ZN(_06588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13637_ (.A1(_06539_),
    .A2(_06549_),
    .ZN(_06589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13638_ (.A1(_06543_),
    .A2(_06548_),
    .B(_06589_),
    .ZN(_06590_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13639_ (.A1(_06586_),
    .A2(_06588_),
    .A3(_06590_),
    .Z(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13640_ (.A1(_06533_),
    .A2(_06550_),
    .Z(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13641_ (.A1(_06533_),
    .A2(_06550_),
    .Z(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13642_ (.A1(_06532_),
    .A2(_06592_),
    .B(_06593_),
    .ZN(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13643_ (.A1(_06536_),
    .A2(_06537_),
    .Z(_06595_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13644_ (.A1(_06536_),
    .A2(_06537_),
    .Z(_06596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13645_ (.A1(_06535_),
    .A2(_06595_),
    .B(_06596_),
    .ZN(_06597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13646_ (.A1(_00387_),
    .A2(_03727_),
    .ZN(_06599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13647_ (.A1(_00397_),
    .A2(_03558_),
    .ZN(_06600_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13648_ (.A1(_06597_),
    .A2(_06599_),
    .A3(_06600_),
    .Z(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13649_ (.A1(_06594_),
    .A2(_06601_),
    .Z(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13650_ (.A1(_06585_),
    .A2(_06591_),
    .A3(_06602_),
    .Z(_06603_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13651_ (.A1(_06581_),
    .A2(_06584_),
    .A3(_06603_),
    .ZN(_06604_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13652_ (.A1(_06575_),
    .A2(_06579_),
    .A3(_06604_),
    .Z(_06605_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13653_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[1] ),
    .A2(_06573_),
    .A3(_06605_),
    .Z(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13654_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[0] ),
    .A2(_06565_),
    .B(_06567_),
    .ZN(_06607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13655_ (.A1(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[0] ),
    .A2(_06565_),
    .ZN(_06608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13656_ (.A1(_06511_),
    .A2(_06607_),
    .B(_06608_),
    .ZN(_06610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13657_ (.A1(_06606_),
    .A2(_06610_),
    .Z(_06611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13658_ (.A1(_05280_),
    .A2(net26),
    .ZN(_06612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13659_ (.A1(_05822_),
    .A2(_06611_),
    .B(_06612_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13660_ (.A1(_05442_),
    .A2(_05387_),
    .B(_00568_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13661_ (.A1(_05463_),
    .A2(_05387_),
    .B(_00570_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13662_ (.A1(_05572_),
    .A2(_05387_),
    .B(_00572_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13663_ (.A1(_06232_),
    .A2(_05387_),
    .B(_00574_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13664_ (.A1(_06146_),
    .A2(_05387_),
    .B(_00576_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13665_ (.D(_00000_),
    .CLK(clknet_leaf_61_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13666_ (.D(_00001_),
    .CLK(clknet_leaf_61_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13667_ (.D(_00002_),
    .CLK(clknet_leaf_62_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13668_ (.D(_00003_),
    .CLK(clknet_leaf_58_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13669_ (.D(_00004_),
    .CLK(clknet_leaf_78_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13670_ (.D(_00005_),
    .CLK(clknet_leaf_78_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13671_ (.D(_00006_),
    .CLK(clknet_leaf_77_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13672_ (.D(_00007_),
    .CLK(clknet_leaf_0_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13673_ (.D(_00008_),
    .CLK(clknet_leaf_0_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13674_ (.D(_00009_),
    .CLK(clknet_leaf_1_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13675_ (.D(_00010_),
    .CLK(clknet_leaf_77_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13676_ (.D(_00011_),
    .CLK(clknet_leaf_3_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13677_ (.D(_00012_),
    .CLK(clknet_leaf_77_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13678_ (.D(_00013_),
    .CLK(clknet_leaf_77_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13679_ (.D(_00014_),
    .CLK(clknet_leaf_0_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13680_ (.D(_00015_),
    .CLK(clknet_leaf_2_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13681_ (.D(_00016_),
    .CLK(clknet_leaf_3_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13682_ (.D(_00017_),
    .CLK(clknet_leaf_0_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13683_ (.D(_00018_),
    .CLK(clknet_leaf_3_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13684_ (.D(_00019_),
    .CLK(clknet_leaf_0_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13685_ (.D(_00020_),
    .CLK(clknet_leaf_0_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13686_ (.D(_00021_),
    .CLK(clknet_leaf_1_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13687_ (.D(_00022_),
    .CLK(clknet_leaf_0_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13688_ (.D(_00023_),
    .CLK(clknet_leaf_2_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13689_ (.D(_00024_),
    .CLK(clknet_leaf_2_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13690_ (.D(_00025_),
    .CLK(clknet_leaf_10_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13691_ (.D(_00026_),
    .CLK(clknet_leaf_8_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13692_ (.D(_00027_),
    .CLK(clknet_leaf_8_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13693_ (.D(_00028_),
    .CLK(clknet_leaf_6_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13694_ (.D(_00029_),
    .CLK(clknet_leaf_6_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13695_ (.D(_00030_),
    .CLK(clknet_leaf_6_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13696_ (.D(_00031_),
    .CLK(clknet_leaf_54_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13697_ (.D(_00032_),
    .CLK(clknet_leaf_57_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13698_ (.D(_00033_),
    .CLK(clknet_leaf_57_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13699_ (.D(_00034_),
    .CLK(clknet_leaf_54_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13700_ (.D(_00035_),
    .CLK(clknet_leaf_64_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13701_ (.D(_00036_),
    .CLK(clknet_leaf_53_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13702_ (.D(_00037_),
    .CLK(clknet_leaf_42_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13703_ (.D(_00038_),
    .CLK(clknet_leaf_47_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13704_ (.D(_00039_),
    .CLK(clknet_leaf_39_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13705_ (.D(_00040_),
    .CLK(clknet_leaf_34_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13706_ (.D(_00041_),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13707_ (.D(_00042_),
    .CLK(clknet_leaf_39_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13708_ (.D(_00043_),
    .CLK(clknet_leaf_33_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13709_ (.D(_00044_),
    .CLK(clknet_leaf_33_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13710_ (.D(_00045_),
    .CLK(clknet_leaf_33_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13711_ (.D(_00046_),
    .CLK(clknet_3_5__leaf_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13712_ (.D(_00047_),
    .CLK(clknet_leaf_13_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13713_ (.D(_00048_),
    .CLK(clknet_leaf_29_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13714_ (.D(_00049_),
    .CLK(clknet_leaf_30_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13715_ (.D(_00050_),
    .CLK(clknet_leaf_14_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13716_ (.D(_00051_),
    .CLK(clknet_leaf_17_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13717_ (.D(_00052_),
    .CLK(clknet_leaf_18_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13718_ (.D(_00053_),
    .CLK(clknet_leaf_21_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13719_ (.D(_00054_),
    .CLK(clknet_leaf_13_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13720_ (.D(_00055_),
    .CLK(clknet_leaf_16_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13721_ (.D(_00056_),
    .CLK(clknet_leaf_20_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13722_ (.D(_00057_),
    .CLK(clknet_leaf_15_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13723_ (.D(_00058_),
    .RN(net36),
    .CLK(clknet_leaf_21_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13724_ (.D(_00059_),
    .RN(net36),
    .CLK(clknet_leaf_36_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13725_ (.D(_00060_),
    .RN(net36),
    .CLK(clknet_leaf_16_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13726_ (.D(_00061_),
    .RN(net36),
    .CLK(clknet_leaf_24_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13727_ (.D(_00062_),
    .RN(net36),
    .CLK(clknet_3_3__leaf_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13728_ (.D(_00063_),
    .RN(net36),
    .CLK(clknet_leaf_37_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13729_ (.D(_00064_),
    .RN(net36),
    .CLK(clknet_leaf_16_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13730_ (.D(_00065_),
    .RN(net36),
    .CLK(clknet_leaf_16_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13731_ (.D(_00066_),
    .RN(net36),
    .CLK(clknet_leaf_17_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13732_ (.D(_00067_),
    .RN(net36),
    .CLK(clknet_leaf_36_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13733_ (.D(_00068_),
    .RN(net36),
    .CLK(clknet_leaf_20_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13734_ (.D(_00069_),
    .RN(net36),
    .CLK(clknet_leaf_23_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13735_ (.D(_00070_),
    .RN(net36),
    .CLK(clknet_leaf_16_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13736_ (.D(_00071_),
    .RN(net36),
    .CLK(clknet_leaf_15_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13737_ (.D(_00072_),
    .RN(net36),
    .CLK(clknet_leaf_13_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13738_ (.D(_00073_),
    .RN(net36),
    .CLK(clknet_leaf_73_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13739_ (.D(_00074_),
    .RN(net36),
    .CLK(clknet_leaf_73_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13740_ (.D(_00075_),
    .RN(net36),
    .CLK(clknet_leaf_69_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13741_ (.D(_00076_),
    .RN(net36),
    .CLK(clknet_leaf_71_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13742_ (.D(_00077_),
    .RN(net36),
    .CLK(clknet_leaf_68_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13743_ (.D(_00078_),
    .RN(net36),
    .CLK(clknet_leaf_68_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13744_ (.D(_00079_),
    .RN(net36),
    .CLK(clknet_leaf_67_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13745_ (.D(_00080_),
    .RN(net36),
    .CLK(clknet_leaf_52_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13746_ (.D(_00081_),
    .RN(net36),
    .CLK(clknet_leaf_51_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13747_ (.D(_00082_),
    .RN(net36),
    .CLK(clknet_leaf_49_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13748_ (.D(_00083_),
    .RN(net36),
    .CLK(clknet_leaf_48_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13749_ (.D(_00084_),
    .RN(net36),
    .CLK(clknet_leaf_48_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13750_ (.D(_00085_),
    .RN(net36),
    .CLK(clknet_leaf_45_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13751_ (.D(_00086_),
    .RN(net36),
    .CLK(clknet_leaf_42_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13752_ (.D(_00087_),
    .RN(net36),
    .CLK(clknet_leaf_43_clk),
    .Q(\DDS_Stage.xPoints_Generator1.CosNew[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13753_ (.D(_00088_),
    .CLK(clknet_leaf_59_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13754_ (.D(_00089_),
    .CLK(clknet_leaf_62_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13755_ (.D(_00090_),
    .CLK(clknet_leaf_59_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13756_ (.D(_00091_),
    .CLK(clknet_leaf_59_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13757_ (.D(_00092_),
    .CLK(clknet_leaf_59_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13758_ (.D(_00093_),
    .CLK(clknet_leaf_58_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13759_ (.D(_00094_),
    .CLK(clknet_leaf_78_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13760_ (.D(_00095_),
    .CLK(clknet_leaf_78_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13761_ (.D(_00096_),
    .CLK(clknet_leaf_78_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13762_ (.D(_00097_),
    .CLK(clknet_leaf_12_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13763_ (.D(_00098_),
    .CLK(clknet_leaf_12_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13764_ (.D(_00099_),
    .CLK(clknet_leaf_1_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _13765_ (.D(_00100_),
    .CLK(clknet_leaf_9_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13766_ (.D(_00101_),
    .CLK(clknet_leaf_10_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13767_ (.D(_00102_),
    .CLK(clknet_leaf_10_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13768_ (.D(_00103_),
    .CLK(clknet_leaf_8_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _13769_ (.D(_00104_),
    .CLK(clknet_leaf_11_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13770_ (.D(_00105_),
    .CLK(clknet_leaf_11_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _13771_ (.D(_00106_),
    .CLK(clknet_leaf_11_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _13772_ (.D(_00107_),
    .CLK(clknet_leaf_10_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13773_ (.D(_00108_),
    .CLK(clknet_leaf_15_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13774_ (.D(_00109_),
    .CLK(clknet_leaf_15_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13775_ (.D(_00110_),
    .CLK(clknet_leaf_6_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13776_ (.D(_00111_),
    .CLK(clknet_leaf_22_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13777_ (.D(_00112_),
    .CLK(clknet_leaf_20_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13778_ (.D(_00113_),
    .CLK(clknet_leaf_15_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13779_ (.D(_00114_),
    .CLK(clknet_leaf_5_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13780_ (.D(_00115_),
    .CLK(clknet_leaf_5_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13781_ (.D(_00116_),
    .CLK(clknet_leaf_4_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13782_ (.D(_00117_),
    .CLK(clknet_leaf_4_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13783_ (.D(_00118_),
    .CLK(clknet_leaf_11_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13784_ (.D(net126),
    .RN(net36),
    .CLK(clknet_leaf_75_clk),
    .Q(\DDS_Stage.LCU.state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13785_ (.D(net130),
    .RN(net36),
    .CLK(clknet_leaf_75_clk),
    .Q(\DDS_Stage.LCU.state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13786_ (.D(_00291_),
    .RN(net36),
    .CLK(clknet_leaf_75_clk),
    .Q(\DDS_Stage.LCU.state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13787_ (.D(\DDS_Stage.LCU.SelMuxConfig ),
    .RN(net36),
    .CLK(clknet_leaf_72_clk),
    .Q(\DDS_Stage.LCU.SelMuxConfigReg ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13788_ (.D(_00119_),
    .RN(net36),
    .CLK(clknet_leaf_63_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13789_ (.D(_00120_),
    .RN(net36),
    .CLK(clknet_leaf_63_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13790_ (.D(_00121_),
    .RN(net36),
    .CLK(clknet_leaf_62_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13791_ (.D(_00122_),
    .RN(net36),
    .CLK(clknet_leaf_73_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13792_ (.D(_00123_),
    .RN(net36),
    .CLK(clknet_leaf_66_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13793_ (.D(_00124_),
    .RN(net36),
    .CLK(clknet_leaf_66_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13794_ (.D(_00125_),
    .RN(net36),
    .CLK(clknet_leaf_65_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13795_ (.D(_00126_),
    .RN(net36),
    .CLK(clknet_leaf_66_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13796_ (.D(_00127_),
    .RN(net36),
    .CLK(clknet_leaf_52_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13797_ (.D(_00128_),
    .RN(net36),
    .CLK(clknet_leaf_50_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13798_ (.D(_00129_),
    .RN(net36),
    .CLK(clknet_leaf_64_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13799_ (.D(_00130_),
    .RN(net36),
    .CLK(clknet_leaf_60_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13800_ (.D(_00131_),
    .RN(net36),
    .CLK(clknet_leaf_60_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13801_ (.D(_00132_),
    .RN(net36),
    .CLK(clknet_leaf_65_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13802_ (.D(_00133_),
    .RN(net36),
    .CLK(clknet_leaf_64_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13803_ (.D(_00134_),
    .RN(net36),
    .CLK(clknet_leaf_63_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13804_ (.D(_00135_),
    .RN(net36),
    .CLK(clknet_leaf_63_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13805_ (.D(_00136_),
    .RN(net36),
    .CLK(clknet_leaf_70_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13806_ (.D(_00137_),
    .RN(net36),
    .CLK(clknet_leaf_73_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13807_ (.D(_00138_),
    .RN(net36),
    .CLK(clknet_leaf_66_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13808_ (.D(_00139_),
    .RN(net36),
    .CLK(clknet_leaf_66_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13809_ (.D(_00140_),
    .RN(net36),
    .CLK(clknet_leaf_66_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13810_ (.D(_00141_),
    .RN(net36),
    .CLK(clknet_leaf_52_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13811_ (.D(_00142_),
    .RN(net36),
    .CLK(clknet_leaf_52_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13812_ (.D(_00143_),
    .RN(net36),
    .CLK(clknet_leaf_50_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13813_ (.D(_00144_),
    .RN(net36),
    .CLK(clknet_leaf_50_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13814_ (.D(_00145_),
    .RN(net36),
    .CLK(clknet_leaf_47_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13815_ (.D(_00146_),
    .RN(net36),
    .CLK(clknet_leaf_46_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13816_ (.D(_00147_),
    .RN(net36),
    .CLK(clknet_leaf_45_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13817_ (.D(_00148_),
    .RN(net36),
    .CLK(clknet_leaf_46_clk),
    .Q(\DDS_Stage.Block_Cosine.agu_1.agu_urgn_in[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13818_ (.D(_00149_),
    .CLK(clknet_leaf_72_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13819_ (.D(_00150_),
    .CLK(clknet_leaf_70_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13820_ (.D(_00151_),
    .CLK(clknet_leaf_71_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13821_ (.D(_00152_),
    .CLK(clknet_leaf_72_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13822_ (.D(_00153_),
    .CLK(clknet_leaf_69_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13823_ (.D(_00154_),
    .CLK(clknet_leaf_68_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13824_ (.D(_00155_),
    .CLK(clknet_leaf_68_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13825_ (.D(_00156_),
    .CLK(clknet_leaf_51_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13826_ (.D(_00157_),
    .CLK(clknet_leaf_51_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13827_ (.D(_00158_),
    .CLK(clknet_leaf_51_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13828_ (.D(_00159_),
    .CLK(clknet_leaf_49_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13829_ (.D(_00160_),
    .CLK(clknet_leaf_48_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13830_ (.D(_00161_),
    .CLK(clknet_leaf_45_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13831_ (.D(_00162_),
    .CLK(clknet_leaf_44_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13832_ (.D(_00163_),
    .CLK(clknet_leaf_43_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegF[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13833_ (.D(_00164_),
    .CLK(clknet_leaf_73_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13834_ (.D(_00165_),
    .CLK(clknet_leaf_70_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13835_ (.D(_00166_),
    .CLK(clknet_leaf_71_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13836_ (.D(_00167_),
    .CLK(clknet_leaf_71_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13837_ (.D(_00168_),
    .CLK(clknet_leaf_68_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13838_ (.D(_00169_),
    .CLK(clknet_leaf_68_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13839_ (.D(_00170_),
    .CLK(clknet_leaf_68_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13840_ (.D(_00171_),
    .CLK(clknet_leaf_51_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13841_ (.D(_00172_),
    .CLK(clknet_leaf_51_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13842_ (.D(_00173_),
    .CLK(clknet_leaf_49_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13843_ (.D(_00174_),
    .CLK(clknet_leaf_49_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13844_ (.D(_00175_),
    .CLK(clknet_leaf_48_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13845_ (.D(_00176_),
    .CLK(clknet_leaf_45_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13846_ (.D(_00177_),
    .CLK(clknet_leaf_42_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _13847_ (.D(_00178_),
    .CLK(clknet_leaf_42_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegP[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13848_ (.D(_00179_),
    .RN(net36),
    .CLK(clknet_leaf_74_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13849_ (.D(_00180_),
    .RN(net36),
    .CLK(clknet_leaf_69_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13850_ (.D(_00181_),
    .RN(net36),
    .CLK(clknet_leaf_71_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13851_ (.D(_00182_),
    .RN(net36),
    .CLK(clknet_leaf_72_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13852_ (.D(_00183_),
    .RN(net36),
    .CLK(clknet_leaf_69_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13853_ (.D(_00184_),
    .RN(net36),
    .CLK(clknet_leaf_67_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13854_ (.D(_00185_),
    .RN(net36),
    .CLK(clknet_leaf_67_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13855_ (.D(_00186_),
    .RN(net36),
    .CLK(clknet_leaf_67_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13856_ (.D(_00187_),
    .RN(net36),
    .CLK(clknet_leaf_51_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13857_ (.D(_00188_),
    .RN(net36),
    .CLK(clknet_leaf_51_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13858_ (.D(_00189_),
    .RN(net36),
    .CLK(clknet_leaf_49_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13859_ (.D(_00190_),
    .RN(net36),
    .CLK(clknet_leaf_48_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13860_ (.D(_00191_),
    .RN(net36),
    .CLK(clknet_leaf_48_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13861_ (.D(_00192_),
    .RN(net36),
    .CLK(clknet_leaf_44_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13862_ (.D(_00193_),
    .RN(net36),
    .CLK(clknet_leaf_42_clk),
    .Q(\DDS_Stage.xPoints_Generator1.RegFrequency[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 _13863_ (.D(_00194_),
    .RN(net36),
    .CLK(clknet_leaf_64_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13864_ (.D(_00195_),
    .RN(net36),
    .CLK(clknet_leaf_63_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13865_ (.D(_00196_),
    .RN(net36),
    .CLK(clknet_leaf_2_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13866_ (.D(_00197_),
    .RN(net36),
    .CLK(clknet_leaf_74_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13867_ (.D(_00198_),
    .RN(net36),
    .CLK(clknet_3_0__leaf_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13868_ (.D(_00199_),
    .RN(net36),
    .CLK(clknet_leaf_65_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13869_ (.D(_00200_),
    .RN(net36),
    .CLK(clknet_leaf_54_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13870_ (.D(_00201_),
    .RN(net36),
    .CLK(clknet_leaf_53_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13871_ (.D(_00202_),
    .RN(net36),
    .CLK(clknet_leaf_52_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13872_ (.D(_00203_),
    .RN(net36),
    .CLK(clknet_leaf_50_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13873_ (.D(_00204_),
    .RN(net36),
    .CLK(clknet_leaf_64_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13874_ (.D(_00205_),
    .RN(net36),
    .CLK(clknet_leaf_60_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 _13875_ (.D(_00206_),
    .RN(net36),
    .CLK(clknet_leaf_55_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13876_ (.D(_00207_),
    .RN(net36),
    .CLK(clknet_leaf_65_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13877_ (.D(_00208_),
    .RN(net36),
    .CLK(clknet_leaf_61_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13878_ (.D(_00209_),
    .RN(net36),
    .CLK(clknet_leaf_63_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13879_ (.D(_00210_),
    .RN(net36),
    .CLK(clknet_leaf_61_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13880_ (.D(_00211_),
    .RN(net36),
    .CLK(clknet_leaf_61_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13881_ (.D(_00212_),
    .RN(net36),
    .CLK(clknet_leaf_62_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13882_ (.D(_00213_),
    .RN(net36),
    .CLK(clknet_leaf_60_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13883_ (.D(_00214_),
    .RN(net36),
    .CLK(clknet_leaf_60_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13884_ (.D(_00215_),
    .RN(net36),
    .CLK(clknet_leaf_59_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13885_ (.D(_00216_),
    .RN(net36),
    .CLK(clknet_leaf_55_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13886_ (.D(_00217_),
    .RN(net36),
    .CLK(clknet_leaf_60_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13887_ (.D(_00218_),
    .RN(net36),
    .CLK(clknet_3_2__leaf_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13888_ (.D(_00219_),
    .RN(net36),
    .CLK(clknet_leaf_37_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13889_ (.D(_00220_),
    .RN(net36),
    .CLK(clknet_leaf_9_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13890_ (.D(_00221_),
    .RN(net36),
    .CLK(clknet_leaf_36_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13891_ (.D(_00222_),
    .RN(net36),
    .CLK(clknet_leaf_11_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13892_ (.D(_00223_),
    .RN(net36),
    .CLK(clknet_leaf_17_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13893_ (.D(_00224_),
    .RN(net36),
    .CLK(clknet_leaf_8_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13894_ (.D(_00225_),
    .RN(net36),
    .CLK(clknet_leaf_17_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13895_ (.D(_00226_),
    .RN(net36),
    .CLK(clknet_leaf_15_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13896_ (.D(_00227_),
    .RN(net36),
    .CLK(clknet_leaf_18_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13897_ (.D(_00228_),
    .RN(net36),
    .CLK(clknet_leaf_15_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13898_ (.D(_00229_),
    .RN(net36),
    .CLK(clknet_leaf_18_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13899_ (.D(_00230_),
    .RN(net36),
    .CLK(clknet_leaf_18_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13900_ (.D(_00231_),
    .RN(net36),
    .CLK(clknet_leaf_19_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13901_ (.D(_00232_),
    .RN(net36),
    .CLK(clknet_leaf_22_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13902_ (.D(_00233_),
    .RN(net36),
    .CLK(clknet_leaf_21_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13903_ (.D(_00234_),
    .RN(net36),
    .CLK(clknet_leaf_20_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13904_ (.D(_00235_),
    .RN(net36),
    .CLK(clknet_leaf_20_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13905_ (.D(_00236_),
    .RN(net36),
    .CLK(clknet_leaf_23_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13906_ (.D(_00237_),
    .RN(net36),
    .CLK(clknet_leaf_23_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13907_ (.D(_00238_),
    .RN(net36),
    .CLK(clknet_leaf_24_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13908_ (.D(_00239_),
    .RN(net36),
    .CLK(clknet_leaf_24_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13909_ (.D(_00240_),
    .RN(net36),
    .CLK(clknet_leaf_24_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13910_ (.D(_00241_),
    .RN(net36),
    .CLK(clknet_leaf_54_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13911_ (.D(_00242_),
    .RN(net36),
    .CLK(clknet_leaf_53_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13912_ (.D(_00243_),
    .RN(net36),
    .CLK(clknet_leaf_54_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13913_ (.D(_00244_),
    .RN(net36),
    .CLK(clknet_leaf_53_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13914_ (.D(_00245_),
    .RN(net36),
    .CLK(clknet_leaf_53_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13915_ (.D(_00246_),
    .RN(net36),
    .CLK(clknet_leaf_53_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13916_ (.D(_00247_),
    .RN(net36),
    .CLK(clknet_leaf_42_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13917_ (.D(_00248_),
    .RN(net36),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13918_ (.D(_00249_),
    .RN(net36),
    .CLK(clknet_leaf_39_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13919_ (.D(_00250_),
    .RN(net36),
    .CLK(clknet_leaf_34_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13920_ (.D(_00251_),
    .RN(net36),
    .CLK(clknet_leaf_32_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13921_ (.D(_00252_),
    .RN(net36),
    .CLK(clknet_leaf_31_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13922_ (.D(_00253_),
    .RN(net36),
    .CLK(clknet_leaf_31_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13923_ (.D(_00254_),
    .RN(net36),
    .CLK(clknet_leaf_33_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13924_ (.D(_00255_),
    .RN(net36),
    .CLK(clknet_leaf_32_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13925_ (.D(_00256_),
    .RN(net36),
    .CLK(clknet_leaf_33_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13926_ (.D(_00257_),
    .RN(net36),
    .CLK(clknet_leaf_28_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13927_ (.D(_00258_),
    .RN(net36),
    .CLK(clknet_leaf_29_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13928_ (.D(_00259_),
    .RN(net36),
    .CLK(clknet_leaf_30_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13929_ (.D(_00260_),
    .RN(net101),
    .CLK(clknet_leaf_28_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13930_ (.D(_00261_),
    .RN(net101),
    .CLK(clknet_leaf_19_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13931_ (.D(_00262_),
    .RN(net101),
    .CLK(clknet_leaf_19_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13932_ (.D(_00263_),
    .RN(net101),
    .CLK(clknet_leaf_19_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13933_ (.D(_00264_),
    .RN(net101),
    .CLK(clknet_leaf_14_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13934_ (.D(_00265_),
    .RN(net101),
    .CLK(clknet_leaf_19_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[-1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13935_ (.D(_00266_),
    .RN(net101),
    .CLK(clknet_leaf_20_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13936_ (.D(_00267_),
    .RN(net101),
    .CLK(clknet_leaf_16_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13937_ (.D(_00268_),
    .RN(net101),
    .CLK(clknet_3_5__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13938_ (.D(_00269_),
    .RN(net101),
    .CLK(clknet_leaf_31_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13939_ (.D(_00270_),
    .RN(net101),
    .CLK(clknet_leaf_31_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13940_ (.D(_00271_),
    .RN(net101),
    .CLK(clknet_leaf_30_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13941_ (.D(_00272_),
    .RN(net101),
    .CLK(clknet_leaf_29_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13942_ (.D(_00273_),
    .RN(net101),
    .CLK(clknet_leaf_29_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13943_ (.D(_00274_),
    .RN(net101),
    .CLK(clknet_leaf_29_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13944_ (.D(_00275_),
    .RN(net101),
    .CLK(clknet_leaf_28_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13945_ (.D(_00276_),
    .RN(net101),
    .CLK(clknet_leaf_27_clk),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13946_ (.D(_00277_),
    .RN(net101),
    .CLK(clknet_3_7__leaf_clk),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13947_ (.D(_00278_),
    .RN(net101),
    .CLK(clknet_leaf_27_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13948_ (.D(_00279_),
    .RN(net101),
    .CLK(clknet_leaf_26_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13949_ (.D(_00280_),
    .RN(net101),
    .CLK(clknet_leaf_26_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13950_ (.D(_00281_),
    .RN(net101),
    .CLK(clknet_leaf_26_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13951_ (.D(_00282_),
    .RN(net101),
    .CLK(clknet_leaf_27_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13952_ (.D(_00283_),
    .RN(net101),
    .CLK(clknet_leaf_26_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13953_ (.D(_00284_),
    .RN(net36),
    .CLK(clknet_leaf_58_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13954_ (.D(_00285_),
    .RN(net36),
    .CLK(clknet_leaf_59_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13955_ (.D(_00286_),
    .RN(net101),
    .CLK(clknet_leaf_56_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _13956_ (.D(_00287_),
    .RN(net101),
    .CLK(clknet_leaf_56_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _13957_ (.D(_00288_),
    .RN(net36),
    .CLK(clknet_leaf_58_clk),
    .Q(\DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clone10 (.I(net88),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 clone11 (.I(net64),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clone12 (.I(net141),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clone13 (.I(net141),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 clone14 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clone18 (.I(net90),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 clone2 (.I(net62),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 clone21 (.I(net78),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clone22 (.I(net146),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clone23 (.I(net146),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 clone31 (.I(net136),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlya_4 clone36 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[15] ),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clone38 (.I(net140),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clone39 (.I(net139),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 clone43 (.I(net144),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 clone44 (.I(net144),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlya_4 clone48 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out[25] ),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 clone5 (.I(_02607_),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlya_4 clone53 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-20] ),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlya_4 clone54 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-20] ),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlya_4 clone56 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-19] ),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlya_4 clone57 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in[-19] ),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clone59 (.I(net159),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 clone6 (.I(net59),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 clone7 (.I(net88),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 clone8 (.I(net76),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 clone9 (.I(net75),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 fanout36 (.I(net19),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold48 (.I(net102),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 hold49 (.I(net19),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(net162),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(FreqPhase[7]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold52 (.I(net14),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(FreqPhase[9]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold54 (.I(net16),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(FreqPhase[8]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold56 (.I(net15),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(FreqPhase[10]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(net3),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(FreqPhase[5]),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold60 (.I(net12),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(FreqPhase[2]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold62 (.I(net9),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(FreqPhase[6]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(net13),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(FreqPhase[4]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold66 (.I(net11),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(net121),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(net10),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(FreqPhase[3]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(net164),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(net163),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(net169),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(_05215_),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(_00289_),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(net166),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(LoadF),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(_05346_),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(_00290_),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(net165),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(net168),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(net167),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(net171),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold83 (.I(rst),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold84 (.I(FreqPhase[13]),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold85 (.I(FreqPhase[0]),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold86 (.I(FreqPhase[1]),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold87 (.I(FreqPhase[11]),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold88 (.I(FreqPhase[14]),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold89 (.I(FreqPhase[12]),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold90 (.I(LoadP),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold91 (.I(_05291_),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold92 (.I(Enable),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1 (.I(net134),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(net119),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(net117),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(net111),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(net115),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(net103),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(net107),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(net105),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(net128),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(net124),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 input19 (.I(net100),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(net122),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(net109),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(net127),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(net132),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(net123),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(net133),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(net131),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(net113),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(Cos_Out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(Cos_Out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(Cos_Out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(Cos_Out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(Cos_Out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(Cos_Out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(Cos_Out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(Cos_Out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(Cos_Out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output29 (.I(net29),
    .Z(Cos_Out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output30 (.I(net30),
    .Z(Cos_Out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output31 (.I(net31),
    .Z(Cos_Out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output32 (.I(net32),
    .Z(Cos_Out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output33 (.I(net33),
    .Z(Cos_Out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output34 (.I(net34),
    .Z(Cos_Out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output35 (.I(net35),
    .Z(Cos_Out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer1 (.I(_02754_),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer10 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-14] ),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 rebuffer11 (.I(_00960_),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 rebuffer12 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-3] ),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer13 (.I(_05149_),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer14 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-14] ),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer15 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-15] ),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer16 (.I(_01076_),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer17 (.I(_03335_),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer18 (.I(_04853_),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer19 (.I(_01095_),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer2 (.I(_04155_),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer20 (.I(_00964_),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer21 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-13] ),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer22 (.I(_00366_),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer23 (.I(_00366_),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 rebuffer24 (.I(_00362_),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer25 (.I(_05740_),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer26 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-13] ),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer27 (.I(_03342_),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer28 (.I(_05083_),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer29 (.I(_05374_),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer3 (.I(_02489_),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer30 (.I(_05133_),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer32 (.I(_00391_),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer33 (.I(net96),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer34 (.I(net96),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer35 (.I(_04859_),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer37 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-3] ),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer4 (.I(_01328_),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer40 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-15] ),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer41 (.I(net139),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer42 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2[-15] ),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 rebuffer45 (.I(_00362_),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlya_1 rebuffer46 (.I(_05445_),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer47 (.I(_00366_),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer49 (.I(_03416_),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer5 (.I(_05199_),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer50 (.I(_02610_),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer51 (.I(_02600_),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer52 (.I(_02597_),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer55 (.I(_01286_),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer58 (.I(_00778_),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer60 (.I(_00366_),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer61 (.I(_01938_),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer62 (.I(net73),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer7 (.I(\DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1[-15] ),
    .Z(net59));
 assign io_oeb[0] = net37;
 assign io_oeb[10] = net47;
 assign io_oeb[11] = net48;
 assign io_oeb[12] = net49;
 assign io_oeb[13] = net50;
 assign io_oeb[14] = net51;
 assign io_oeb[15] = net52;
 assign io_oeb[1] = net38;
 assign io_oeb[2] = net39;
 assign io_oeb[3] = net40;
 assign io_oeb[4] = net41;
 assign io_oeb[5] = net42;
 assign io_oeb[6] = net43;
 assign io_oeb[7] = net44;
 assign io_oeb[8] = net45;
 assign io_oeb[9] = net46;
endmodule

