* NGSPICE file created from DDS_Module.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_16 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_20 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_1 I Z VDD VNW VPW VSS
.ends

.subckt DDS_Module Cos_Out[0] Cos_Out[10] Cos_Out[11] Cos_Out[12] Cos_Out[13] Cos_Out[14]
+ Cos_Out[15] Cos_Out[1] Cos_Out[2] Cos_Out[3] Cos_Out[4] Cos_Out[5] Cos_Out[6] Cos_Out[7]
+ Cos_Out[8] Cos_Out[9] Enable FreqPhase[0] FreqPhase[10] FreqPhase[11] FreqPhase[12]
+ FreqPhase[13] FreqPhase[14] FreqPhase[15] FreqPhase[1] FreqPhase[2] FreqPhase[3]
+ FreqPhase[4] FreqPhase[5] FreqPhase[6] FreqPhase[7] FreqPhase[8] FreqPhase[9] LoadF
+ LoadP clk io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[15] io_oeb[1] io_oeb[2]
+ io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] rst vdd vss
+ io_oeb[14] io_oeb[13]
XFILLER_0_20_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06883_ _05420_ _05680_ _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09671_ _02553_ _02557_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07534__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08622_ _00428_ _01508_ _01520_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_49_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08553_ _01389_ _01417_ _01451_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09287__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07504_ _05431_ _06779_ _00455_ _05658_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11094__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08484_ _00385_ net156 _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11094__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07837__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07435_ _05409_ _05420_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09039__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07366_ _00403_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09105_ _00373_ _06672_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07297_ _05387_ _00346_ _00349_ _00350_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_131_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09036_ _01852_ _01928_ _01929_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07494__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09762__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07507__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09938_ _02772_ _02821_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09869_ _02749_ _02753_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07525__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11900_ _00387_ _01956_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12880_ _00365_ _03558_ _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11831_ _04651_ _04672_ _04673_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09278__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07828__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11762_ _04601_ _04603_ _04604_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_36_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11624__A3 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13501_ _05822_ _06441_ _06442_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10713_ _03501_ _03504_ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11693_ _04534_ _04535_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13432_ _06367_ _06368_ _06369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_10644_ _00388_ _00385_ _06744_ _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11388__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10575_ _03389_ _03390_ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13363_ _06216_ _06294_ _06295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xrebuffer7 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-15\] net59 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07300__I1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12314_ _05146_ _05156_ _05157_ _05158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_23_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13294_ _06143_ _06219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_146_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12245_ _05074_ _05077_ _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12176_ _04397_ _04398_ _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10899__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11560__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11127_ _03915_ _03968_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11058_ _00365_ _03018_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12104__A4 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10009_ _02808_ _02818_ _02891_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_87_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10823__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07579__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07220_ _05409_ _06614_ _05658_ _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_116_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07151_ _06232_ _06734_ _06768_ _06769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_3_2__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07082_ _05822_ _06708_ _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12879__A2 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11000__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09744__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11551__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07984_ _00883_ _00884_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09723_ _00355_ _06742_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06935_ _06232_ _05875_ _06243_ _06254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__12500__A1 _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ _02459_ _02463_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06866_ _05420_ _05496_ _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_97_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08605_ _01450_ _01452_ _01503_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_49_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09585_ _02372_ _02373_ _02472_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08536_ _00424_ _01433_ _01434_ _01426_ _01317_ _00418_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_4
XFILLER_0_77_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10409__A4 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08467_ _01262_ _01266_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10908__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08483__A2 _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11082__A4 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07418_ _06232_ _06621_ _06676_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08398_ _01276_ _01298_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_52_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07349_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-3\] _00390_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_116_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10360_ _03196_ _03238_ _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07994__A1 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09019_ _01842_ _01858_ _01912_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10291_ _03085_ _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_20_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12030_ _00387_ _01794_ _04873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_148_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12932_ _05823_ _05828_ _05829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_137_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08171__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12863_ _05692_ _05716_ _05752_ _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11058__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11814_ net70 _01430_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12794_ _05571_ _05573_ _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_139_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10805__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11745_ _04579_ _04587_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08474__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11676_ _04518_ _04512_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12558__A1 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13415_ _06347_ _06348_ _06349_ _06350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_40_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10627_ _00398_ _06730_ _06738_ _00394_ _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_36_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08226__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13346_ _00381_ _03558_ _06277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10558_ net63 _06730_ net57 _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_134_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13277_ _06041_ _06108_ _06202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10489_ net57 _02704_ _03365_ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_59_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12228_ _04365_ _04369_ _05070_ _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12159_ _04999_ _05000_ _05002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_120_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11049__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11049__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _00379_ _06674_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12797__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08321_ _01222_ _01221_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08252_ _01147_ _01148_ _01153_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_7_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07203_ _05420_ _05550_ _06774_ _06813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12549__A1 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _01024_ _01063_ _01084_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07134_ _05572_ _06092_ _06753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_43_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11772__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07065_ _05409_ _05594_ _06693_ _06694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09717__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10327__A3 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11524__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12721__A1 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07772__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07967_ _00769_ _00867_ _00868_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_156_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06951__A2 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ _02513_ _02510_ _02539_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06918_ _05442_ _05452_ _06070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07898_ _00785_ _00798_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08153__A1 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08153__B2 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09637_ _02519_ _02523_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06849_ DDS_Stage.LCU.state\[1\] _05160_ _05324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07504__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09568_ _02452_ _02455_ _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_26_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12788__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _01366_ _01418_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_148_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09499_ _02338_ _02387_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_148_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11530_ _04314_ _04315_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11460__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11461_ _00361_ _02236_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09405__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_122_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__B2 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13200_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-6\] _06118_ _06119_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_10412_ _03209_ _03289_ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_135_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10015__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11392_ _04195_ _04196_ _04197_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_150_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13131_ _05985_ _06000_ _06044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10343_ _00379_ _06742_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13062_ _03485_ _00378_ _05969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10274_ _03112_ _03153_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11515__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12013_ _04147_ _04160_ _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07195__A2 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_131_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11279__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12915_ _03018_ _00387_ _05810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09892__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08695__A2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07498__A3 _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13895_ _00226_ net36 clknet_leaf_15_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09892__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12846_ _05447_ _05537_ _05733_ _05735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_TAPCELL_ROW_83_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12777_ _05659_ _05568_ _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_140_Left_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11451__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11728_ _04556_ _04559_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11451__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11659_ _04441_ _04454_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11203__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13329_ _06186_ _06257_ _06258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11506__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ _01740_ _01765_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08383__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07186__A2 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07821_ _06059_ _00569_ _00726_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07752_ net104 DDS_Stage.xPoints_Generator1.RegP\[-8\] _00684_ _00692_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07683_ DDS_Stage.xPoints_Generator1.RegFrequency\[-4\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-4\]
+ _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_125_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08686__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09422_ _02155_ _02139_ _02225_ _02311_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__10493__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09353_ _02170_ _02222_ _02242_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09635__A1 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08304_ _01205_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10245__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09284_ _02105_ _02108_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08235_ _01098_ _01122_ _01136_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_145_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08166_ _01038_ _01066_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12942__A1 _05336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07117_ _06059_ _06737_ _06739_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08097_ net61 _05833_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_37_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07048_ _05822_ _06679_ _06680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10921__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08999_ _01822_ _01830_ _01892_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06924__A2 _06125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09469__A4 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10961_ _03802_ _03803_ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07234__C _06006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08677__A2 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12700_ _05494_ _05495_ _05577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_70_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13680_ _00015_ clknet_leaf_2_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10892_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-24\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-24\]
+ _05171_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12631_ _05467_ _05501_ _05502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10236__A2 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12562_ _05411_ _05426_ _05427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_148_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11513_ _04296_ _04300_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12493_ _05353_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11444_ _04251_ _04252_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_22_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09929__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11197__B1 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11375_ _04215_ _04216_ _04217_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13114_ _06021_ _06022_ _06025_ _06026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_10326_ net63 _06708_ net57 _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07409__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13045_ _05881_ _05895_ _05950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10257_ _03135_ _03136_ _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07168__A2 _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10188_ _03060_ _03068_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09314__B1 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13947_ _00278_ net101 clknet_leaf_27_clk net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08668__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13661__A2 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11672__A1 _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13878_ _00209_ net36 clknet_leaf_63_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_72_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06983__C _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12829_ _05692_ _05716_ _05717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13413__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11424__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09093__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11975__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08020_ _00918_ _00921_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_53_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06851__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08053__B1 _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09971_ _05280_ _02854_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08922_ _01741_ _01815_ _01816_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12152__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08853_ _01673_ _01677_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10163__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06906__A2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07804_ net60 DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[19\] _00395_ _00718_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08784_ _01656_ _01680_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08108__A1 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07735_ _00682_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_123_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08659__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10466__A2 _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07666_ DDS_Stage.xPoints_Generator1.CosNew\[-6\] _00633_ _00577_ _00634_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09405_ _06642_ _00398_ _00394_ _06649_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13892__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13404__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07597_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[30\] _00575_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11415__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09336_ _02225_ _02226_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__12612__B1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11966__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07095__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09267_ _02065_ _02132_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_138_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06842__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08218_ _01038_ _01066_ _00986_ _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_50_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09198_ _02006_ _02088_ _02089_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12915__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11718__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ _00355_ _06598_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07398__A2 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11160_ _03933_ _04001_ _04002_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10111_ _02895_ _02910_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09139__A3 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11091_ _00361_ _03266_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10042_ _02856_ _02857_ _02923_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__10154__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold52 net14 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold63 FreqPhase[6] net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold74 _00289_ net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold85 FreqPhase[0] net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_98_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13801_ _00132_ net36 clknet_leaf_65_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11993_ _04123_ _04125_ _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09847__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13732_ _00067_ net36 clknet_leaf_36_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_10944_ _03788_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13883__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13663_ _06232_ _05387_ _00574_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10875_ _03031_ _03637_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12614_ _05479_ _05482_ _05483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13594_ _06542_ _06543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_14_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12545_ _04022_ _04030_ _05407_ _05408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12476_ _05298_ _05327_ _05332_ _05334_ _05336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_124_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11427_ _04256_ _04269_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_78_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11358_ _00375_ _01693_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10309_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[22\] _03189_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11289_ _04129_ _04130_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13028_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-8\] _05932_ _05933_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07010__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07561__A2 _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer17 _03335_ net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer28 _05083_ net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09838__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07520_ _05182_ _00520_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13874__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07451_ _05518_ _05789_ _06070_ _06721_ _05658_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_88_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07382_ _00411_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_146_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09121_ _01923_ _01936_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07077__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09052_ _01801_ _01944_ _01945_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_100_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08003_ _00904_ _00890_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09954_ _02834_ _02837_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13322__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12125__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08905_ _01712_ _01713_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09885_ _02767_ _02768_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07001__A1 _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08836_ _06633_ _00385_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07780__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08767_ _01578_ _01663_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_79_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07718_ net116 DDS_Stage.xPoints_Generator1.RegF\[-9\] _00667_ _00674_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08698_ _01587_ _01595_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13865__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07649_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-9\] DDS_Stage.xPoints_Generator1.RegFrequency\[-9\]
+ _00614_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07512__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07855__A3 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13389__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10660_ _03529_ _03534_ _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_137_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07068__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09319_ net60 _06696_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10591_ _03422_ _03466_ _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08624__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12330_ _05175_ _05176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_23_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12261_ _05101_ _05102_ _05103_ _05104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08568__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11212_ _04052_ _04054_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_32_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12192_ _04379_ _04380_ _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput20 net20 Cos_Out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput31 net31 Cos_Out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07240__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11143_ net86 _03485_ _03416_ net84 _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13313__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11074_ _03898_ _03911_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10025_ _02902_ _02906_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07543__A2 _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11976_ _04816_ _04817_ _04818_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_85_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09296__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13856__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13715_ _00050_ clknet_leaf_14_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10927_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-8\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-8\]
+ _05171_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13646_ _00387_ _03727_ _06599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10858_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[5\] _03728_ _03729_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_30_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12052__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13577_ _06473_ _06477_ _06525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10789_ _03589_ _03592_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_147_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12528_ _05384_ _05389_ _05390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_136_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12459_ _05016_ _05316_ _05317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09220__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07231__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12107__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ _05822_ net152 _06427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11866__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09670_ _02554_ _02555_ _02556_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06882_ _05550_ _05669_ _05680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_118_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07534__A2 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08621_ _01510_ _01519_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08552_ _01392_ _01416_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09287__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07503_ _05409_ _05995_ _06761_ _06146_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08483_ _00388_ _06416_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11094__A2 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07434_ _05658_ _06830_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09039__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07365_ DDS_Stage.xPoints_Generator1.CosNew\[-15\] DDS_Stage.xPoints_Generator1.RegP\[-15\]
+ _00402_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone11_I net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08798__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09104_ _01995_ _01996_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07296_ _05658_ _06687_ _05171_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09035_ net61 net60 _06672_ _06674_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07470__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07222__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09937_ _02799_ _02820_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07507__C _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09868_ _02591_ _02750_ _02751_ _02752_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__07525__A2 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08819_ _01656_ _01680_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09799_ _02650_ _02651_ _02683_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11830_ _04670_ _04671_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09278__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11761_ _04484_ _04503_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07242__C _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13500_ _05280_ net23 _06442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11624__A4 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10712_ _03311_ _03525_ _03585_ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11692_ _04525_ _04530_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13431_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-4\] _06293_ _06215_ _06368_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10643_ _03516_ _03517_ _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13362_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-4\] _06293_ _06294_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10574_ _03389_ _03390_ _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_134_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12313_ _05154_ _05155_ _05157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13293_ _06132_ _06199_ _06218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_58_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12244_ _05084_ _05085_ _05086_ _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07213__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12175_ _04397_ _04398_ _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10899__A2 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-21\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07213__B2 _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11126_ _03915_ _03968_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11057_ _00361_ _03189_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08713__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10008_ _02811_ _02815_ _02816_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_64_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11959_ _04759_ _04792_ _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_87_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13629_ _00387_ _03725_ _06545_ _06580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_17_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _06243_ _06469_ _06146_ _06768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_82_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07452__A1 _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07081_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-1\] _06708_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09874__I _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07204__A1 _06646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11000__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08952__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07983_ _00883_ _00884_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09722_ _02607_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06934_ _05572_ _05886_ _06243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11839__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09823__B _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09653_ _02514_ _02539_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06865_ _05474_ _05485_ _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__10511__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08604_ _01474_ _01502_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clone59_I net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09584_ _00373_ _06691_ _02374_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08535_ _01349_ _01425_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_148_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08466_ _01364_ _01299_ _01365_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07417_ _06059_ _00435_ _00436_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08397_ _01278_ _01291_ _01297_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_80_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07348_ _00389_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_21_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10578__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07443__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07279_ _05822_ _00331_ _00334_ _00335_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07994__A2 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09018_ _01844_ _01857_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10290_ _03166_ _03169_ _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10750__A1 _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09499__A2 _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12931_ _05825_ _05827_ _05828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08171__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12862_ _05657_ _05690_ _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11813_ _04647_ _04655_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11058__A2 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12793_ _03189_ _00378_ _05586_ _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_29_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11744_ _04580_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11675_ _04508_ _04517_ _04507_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_81_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13414_ _00381_ _03679_ _06349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12558__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10626_ _02704_ _03499_ _03500_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_40_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13345_ _03556_ _00384_ _06275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07434__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ net63 _06730_ net57 _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13276_ _06043_ _06107_ _06201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10488_ net63 _06730_ _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12227_ _04360_ _04364_ _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12158_ _04999_ _05000_ _05001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11109_ _03885_ _03895_ _03951_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12089_ _04930_ _04931_ _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_75_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08259__B _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11049__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08320_ _00947_ _00973_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12797__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08251_ _01149_ _01150_ _01152_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ _05518_ _06340_ _06721_ _05778_ _05658_ _06812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__12549__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08182_ _01049_ _01062_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07133_ _06751_ _06752_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07425__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11772__A3 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07064_ _05420_ _06681_ _06693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10980__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08925__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12721__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07966_ _00822_ _00866_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09705_ _02562_ _02569_ _02590_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06917_ _05280_ _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
X_07897_ _00785_ _00798_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08153__A2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09636_ _02520_ _02521_ _02522_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06848_ _05280_ _05302_ _05193_ _05237_ _05313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_136_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12237__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09567_ _02453_ _02454_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_26_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12788__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08518_ _01389_ _01417_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09498_ _02365_ _02386_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08449_ _01348_ _01328_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_148_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11460__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11460_ _00365_ _02153_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09405__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10411_ _03285_ _03288_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07416__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11391_ _04229_ _04233_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_116_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13130_ _05946_ _06003_ _06042_ _06043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10342_ _03219_ _03220_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13061_ _05870_ _05966_ _05967_ _05968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10273_ _03131_ _03152_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12012_ _04838_ _04842_ _04854_ _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11279__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09341__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12914_ _05709_ _05807_ _05808_ _05809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13894_ _00225_ net36 clknet_leaf_17_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_88_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12845_ _05632_ _05727_ _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_83_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12776_ _05565_ _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11727_ _04567_ _04568_ _04569_ _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11451__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11658_ _04498_ _04499_ _04500_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_126_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10609_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[26\] _03485_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_4_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11203__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11589_ _04190_ _04191_ _04189_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_52_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13328_ _06191_ _06257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08080__A1 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13259_ _06178_ _06182_ _06183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_110_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07820_ _05280_ _00388_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08383__A2 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07751_ _00691_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07682_ _00647_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09421_ _02157_ _02158_ _02224_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__10493__A3 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09352_ _02172_ _02221_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09635__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08303_ _01200_ _01203_ _01204_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_19_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09283_ _02087_ _02095_ _02173_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_145_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08234_ _01133_ _01135_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08165_ _01038_ _01066_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07249__I1 _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07116_ _05822_ _06738_ _06739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08096_ _00363_ _05864_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10953__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07047_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-6\] _06679_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09020__B1 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10705__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08998_ _01825_ _01829_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07949_ _00807_ _00849_ _00850_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_67_clk clknet_3_1__leaf_clk clknet_leaf_67_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09323__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10960_ _00381_ net135 _02499_ _00384_ _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11130__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08677__A3 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09619_ _02474_ _02475_ _02505_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10891_ _03760_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12630_ _05486_ _05500_ _05501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_65_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07531__B _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12561_ _05416_ _05425_ _05426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_148_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11512_ _04321_ _04341_ _04354_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_156_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12492_ net20 _05352_ _05171_ _05353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_156_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11443_ _04187_ _04221_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_110_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09929__A3 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11197__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11197__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11374_ _00387_ _01430_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13113_ _05927_ _06024_ _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10325_ _03200_ _03203_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13044_ _05869_ _05880_ _05949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10256_ _02966_ _03046_ _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ _03063_ _03067_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12449__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-24\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07425__C _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_clk clknet_3_3__leaf_clk clknet_leaf_58_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09314__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09314__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13946_ _00277_ net101 clknet_3_7__leaf_clk net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_88_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13877_ _00208_ net36 clknet_leaf_61_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XANTENNA__07441__B _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12828_ _05695_ _05699_ _05715_ _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__06836__I _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11424__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12759_ _05543_ _05640_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_96_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08053__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08053__B2 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09970_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[18\] _02854_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_0_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08921_ _01744_ _01747_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08852_ _01741_ _01744_ _01747_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_127_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11360__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10163__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07803_ _05387_ _00358_ _00717_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08783_ _01664_ _01666_ _01679_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08108__A2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_49_clk clknet_3_1__leaf_clk clknet_leaf_49_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07734_ net7 DDS_Stage.xPoints_Generator1.RegF\[-1\] _00667_ _00682_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_140_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07665_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-6\] DDS_Stage.xPoints_Generator1.RegFrequency\[-6\]
+ _00632_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09404_ _02213_ _02292_ _02293_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_9_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07596_ _05387_ _00573_ _00574_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_105_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09335_ _02157_ _02158_ _02224_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__12612__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11415__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12612__B2 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07778__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09266_ _02068_ _02131_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07095__A2 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08217_ _01097_ _01117_ _01118_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_106_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09197_ _02007_ _02008_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_133_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12915__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08148_ net137 _06618_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08079_ _00930_ _00980_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_140_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10110_ _02947_ _02991_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11090_ _00369_ _03018_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09139__A4 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09544__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ _02856_ _02857_ _02923_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10154__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold53 FreqPhase[9] net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold64 net13 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold75 net166 net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold86 FreqPhase[1] net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_13800_ _00131_ net36 clknet_leaf_60_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11992_ _04816_ _04833_ _04834_ _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09847__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13731_ _00066_ net36 clknet_leaf_17_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10943_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[0\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[0\]
+ _05171_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_63_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10874_ _03401_ _03694_ _03744_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13662_ _05572_ _05387_ _00572_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12613_ _05480_ _05481_ _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13593_ _06540_ _06495_ _06541_ _06542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12603__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07688__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12544_ _04025_ _05406_ _05407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12475_ _05285_ _05286_ _05333_ _05328_ _05334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_53_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11426_ _04264_ _04268_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_78_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11357_ _04195_ _04198_ _04199_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_120_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12119__B1 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10308_ _03184_ _03187_ _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_91_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11288_ _04129_ _04130_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_91_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13027_ _05928_ _05931_ _05932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10239_ _02608_ _02704_ _03118_ _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_83_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_21_clk_I clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer18 _04853_ net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_16_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer29 _05374_ net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__09838__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07849__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12842__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13929_ _00260_ net101 clknet_leaf_28_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_77_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08510__A2 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07450_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-15\] _00463_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_36_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07381_ DDS_Stage.xPoints_Generator1.CosNew\[-7\] DDS_Stage.xPoints_Generator1.RegP\[-7\]
+ _00402_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_33_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09120_ _01994_ _02012_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_128_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08274__A1 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07077__A2 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10081__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09051_ _01803_ _01862_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_100_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08002_ _00903_ _00898_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09953_ _02835_ _02836_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_110_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13322__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08904_ _01709_ _01710_ _01708_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11333__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09884_ _02738_ _02746_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07001__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08835_ _06627_ _00388_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13086__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08766_ _01659_ _01662_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07717_ _00673_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08697_ _01590_ _01594_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_68_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07648_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-9\] DDS_Stage.xPoints_Generator1.RegFrequency\[-9\]
+ _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07855__A4 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13389__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07579_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[23\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-8\]
+ _00395_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10927__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09318_ net91 _06691_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07068__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10590_ _03460_ _03465_ _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_11_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10072__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09249_ net56 _01348_ _01700_ _02053_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12260_ _05087_ _05100_ _05103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08017__A1 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11211_ _00372_ _02586_ _02584_ _00375_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08568__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09765__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12191_ _05026_ _05031_ _05033_ _05034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11572__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 net21 Cos_Out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput32 net32 Cos_Out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11142_ _03936_ _03944_ _03984_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07240__A2 _06698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13313__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11073_ _03898_ _03911_ _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10024_ _02902_ _02906_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13077__A1 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12824__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11975_ _00365_ _02586_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13714_ _00049_ clknet_leaf_30_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10926_ _03779_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13937__CLK clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10857_ _03683_ _03719_ _03717_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13645_ _06535_ _06595_ _06596_ _06597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_156_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09697__I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08256__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10788_ _03634_ _03660_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13576_ _06522_ _06524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12052__A2 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12527_ _05385_ _05386_ _05388_ _05389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_26_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08008__A1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12458_ _05287_ _05229_ _05234_ _05316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11409_ _04194_ _04206_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12389_ _05017_ _05234_ _05240_ _05241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_78_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07231__A2 _06125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13792__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12107__A3 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06950_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-20\] _06416_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_20_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06990__A1 _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06881_ _05442_ _05463_ _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__11866__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08620_ _01513_ _01518_ _01425_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08551_ _01448_ _01449_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__12815__A1 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07502_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-6\] _00506_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08482_ _00382_ _06598_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07433_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-18\] _00449_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_102_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10747__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08247__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07364_ _00401_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13240__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_99_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09103_ _01840_ _01920_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10054__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09995__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07295_ _06491_ _00347_ _00348_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_115_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09034_ net61 _06672_ _06674_ net60 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11554__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09936_ _02801_ _02803_ _02819_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__11306__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06981__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09867_ _02589_ _02653_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08818_ _01712_ _01713_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_146_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09798_ _02682_ _02649_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08749_ _06633_ _00382_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11760_ _04592_ _04596_ _04602_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10711_ _00382_ _03520_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_138_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11691_ _04533_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10642_ _03373_ _03440_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13430_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-4\] _06293_ _06367_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_125_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13361_ _06290_ _06292_ _06293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10573_ _03447_ _03448_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12312_ _05154_ _05155_ _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13292_ _06134_ _06198_ _06217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12243_ _05071_ net80 _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12174_ _04943_ _05016_ _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__07213__A2 _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10405__B net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11125_ _03948_ _03967_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11056_ _00369_ _02940_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08713__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10007_ _02867_ _02889_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_87_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11958_ _04794_ _04797_ _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10909_ _03770_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11889_ _04644_ _04675_ _04697_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_73_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13628_ _06533_ _06578_ _06579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06844__I _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13559_ _06459_ _06505_ _06506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11784__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07080_ _05658_ _06706_ _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11536__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08401__A1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08952__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07982_ _00398_ _05398_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06963__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09721_ _00352_ _06744_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_38_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06933_ _05409_ _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_16
XANTENNA__11839__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09901__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06864_ _05431_ _05452_ _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09652_ _02530_ _02538_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10511__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08603_ _01477_ _01501_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09583_ _02367_ _02385_ _02470_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08534_ net56 _01348_ _01432_ _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08465_ _01276_ _01298_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07140__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07416_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-22\] _00436_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08396_ _00885_ _01296_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09968__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07347_ _00387_ _00388_ _05182_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_21_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10578__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11775__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07786__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07278_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-2\] _00335_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09017_ _01893_ _01896_ _01910_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_60_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07518__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06954__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09919_ _02617_ _02714_ _02802_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07534__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12930_ _05641_ _05826_ _05827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12861_ _05747_ _05750_ _05751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_29_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11812_ _04646_ _04648_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08459__A1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12792_ _05584_ _05585_ _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10266__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11743_ _04540_ _04584_ _04585_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07131__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11674_ _04505_ _04506_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_81_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13413_ _00384_ _03558_ _06348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10625_ net63 _06738_ net57 _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_24_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10556_ _03428_ _03431_ _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13344_ _03485_ _00387_ _06274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10487_ _03115_ _03363_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13275_ _06132_ _06199_ _06200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11518__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12226_ _05063_ _05066_ _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_121_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13747__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12157_ _04916_ _04924_ _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_9_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06945__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11108_ _03888_ _03894_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12088_ _04803_ _04828_ _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_88_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11039_ _03854_ _03880_ _03881_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08259__C _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09647__B1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07122__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08250_ net58 _05864_ _01151_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_117_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07201_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-15\] _06811_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_89_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08181_ _01077_ _01082_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_144_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07132_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-25\] _06752_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08622__A1 _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07425__A2 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07063_ _06059_ _06690_ _06692_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11772__A4 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10980__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13738__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_151_Right_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08925__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07965_ _00822_ _00866_ _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09704_ _02512_ _02561_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06916_ _06039_ _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07896_ _00789_ _00797_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10496__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09635_ net143 _06724_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06847_ net18 _05302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13910__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12237__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09566_ _00376_ _06691_ _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08517_ _01392_ _01416_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_77_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07113__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09497_ _02367_ _02385_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_66_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08448_ _01334_ _01337_ _01347_ _01324_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_92_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ net91 net143 _06637_ _06633_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_74_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10935__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10410_ _03286_ _03287_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11390_ _04230_ _04231_ _04232_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_60_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ _03044_ _03128_ _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13060_ _05871_ _05872_ _05967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_60_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10272_ _03134_ _03137_ _03151_ _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__13729__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12011_ _04840_ _04841_ _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_103_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11279__A3 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10487__A1 _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12913_ _05710_ _05711_ _05808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_88_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13893_ _00224_ net36 clknet_leaf_8_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_69_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13901__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12844_ _05822_ net31 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10239__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12775_ _05655_ _05656_ _05657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07104__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11726_ _04553_ _04566_ _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11657_ _04496_ _04497_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_126_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _03481_ _03483_ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11588_ _04426_ _04429_ _04430_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13327_ _06236_ _06255_ _06256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08080__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10539_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[25\] _03416_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_122_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13258_ _06180_ _06181_ _06182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07158__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12209_ _00381_ _00384_ _01956_ _01794_ _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_110_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06918__A1 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13189_ _06106_ _06107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11911__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07750_ net116 DDS_Stage.xPoints_Generator1.RegP\[-9\] _00684_ _00691_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13664__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07681_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-4\] _00646_ _00395_ _00647_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09420_ _02306_ _02309_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_149_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09351_ _02168_ _02169_ _02240_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09096__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11978__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08302_ net155 _00370_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09282_ _02090_ _02094_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08233_ _01134_ _01110_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08164_ _01043_ _01065_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_145_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10402__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07115_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[3\] _06738_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_141_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08095_ _00357_ _06179_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10953__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07046_ _05658_ _06677_ _06678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09020__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09020__B2 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06909__A1 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10705__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11902__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08997_ _01832_ _01860_ _01890_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ net92 net142 _06627_ _06618_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09323__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07879_ _00363_ _06598_ _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11130__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08677__A4 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09618_ _02504_ _02473_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10890_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-25\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-25\]
+ _05171_ _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07304__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09549_ _02423_ _02436_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08834__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12560_ _05419_ _05424_ _05425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11511_ _04290_ _04353_ _04320_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_156_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12491_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-14\] _05279_ _05351_ _05352_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_156_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11442_ _04254_ _04284_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09929__A4 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11197__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11373_ _00381_ _01610_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10324_ _03037_ _03202_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13112_ _06023_ _05926_ _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13043_ _05898_ _05921_ _05947_ _05948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10255_ _03042_ _03045_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09011__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10186_ _03064_ _03065_ _03066_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__13646__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09314__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13945_ _00276_ net101 clknet_leaf_27_clk net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_88_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13876_ _00207_ net36 clknet_leaf_65_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_72_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12827_ _05705_ _05714_ _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12758_ _05387_ _05638_ _05639_ _05640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_127_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10632__A1 _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11709_ _04544_ _04548_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12689_ _00359_ _03558_ _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08053__A2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07169__B _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08920_ _01744_ _01747_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08851_ _01745_ _01746_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_71_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_127_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10163__A3 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11360__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07802_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[18\] _00717_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08782_ _01670_ _01678_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07733_ _00681_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07664_ _00630_ _00631_ _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09403_ _06649_ net58 net95 _06710_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_138_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07595_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-2\] _05182_ _00574_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09334_ _02157_ _02158_ _02224_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__12612__A2 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11415__A3 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09265_ _02155_ _02139_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08216_ _01115_ _01116_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_138_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09196_ _02007_ _02008_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_117_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08147_ _01025_ _01033_ _01048_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07794__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07252__B1 _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08078_ _00945_ _00978_ _00979_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_30_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07029_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-9\] _06664_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10040_ _02860_ _02863_ _02922_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09544__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07526__C _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07555__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold54 net16 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold65 FreqPhase[4] net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold76 LoadF net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold87 FreqPhase[11] net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_11991_ _04817_ _04818_ _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_98_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08504__B1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13730_ _00065_ net36 clknet_leaf_16_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10942_ _03787_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10862__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13661_ _05463_ _05387_ _00570_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_119_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10873_ _03082_ _03695_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12612_ _03485_ _00361_ _00365_ net148 _05481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_149_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13592_ _06493_ _06494_ _06541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12603__A2 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12543_ _04029_ _05406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12474_ _05222_ _05228_ _05333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11425_ _04265_ _04266_ _04267_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_105_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_128_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11356_ _04196_ _04197_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12119__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12119__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10307_ _03186_ _03104_ _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_91_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11287_ _00365_ _02762_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_91_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07209__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13026_ _05829_ _05840_ _05929_ _05931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10238_ net63 _06708_ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07546__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10169_ _02987_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_109_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer19 _01095_ net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13928_ _00259_ net36 clknet_leaf_30_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_137_Left_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07849__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13859_ _00190_ net36 clknet_leaf_48_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_53_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07380_ _00410_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10605__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08274__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09471__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09050_ _01803_ _01862_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10081__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08001_ _00899_ _00902_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09952_ _02684_ _02748_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08903_ _01797_ _01775_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09883_ _02690_ _02737_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11333__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07537__B2 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08834_ _06637_ _00382_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08765_ _01660_ _01661_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13086__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07716_ net112 DDS_Stage.xPoints_Generator1.RegF\[-10\] _00667_ _00673_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11097__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08696_ _01591_ _01592_ _01593_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_95_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07647_ _00617_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13389__A3 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ _00563_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09317_ _00357_ _06701_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09462__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_153_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10072__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09248_ _02138_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_145_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08017__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09214__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09179_ _00373_ _06672_ _02001_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10943__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11210_ _00378_ _02499_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12190_ _05020_ _05032_ _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09765__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12443__B DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-25\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 Cos_Out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__11572__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput33 net33 Cos_Out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11141_ _03939_ _03943_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11072_ _03853_ _03913_ _03914_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07528__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12521__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10023_ _02903_ _02904_ _02905_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__13077__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11974_ _00361_ _02762_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10135__I0 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12824__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10835__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13713_ _00048_ clknet_leaf_29_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10925_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-9\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-9\]
+ _05171_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13644_ _06536_ _06537_ _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_116_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10856_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[31\] _03727_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13575_ _06520_ _06521_ _06522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08256__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10787_ _03652_ _03659_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_125_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12526_ net148 _00361_ _05388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12457_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-21\] _05292_ _05307_ _05312_
+ _05314_ _05315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__08008__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11408_ _04237_ _04250_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12388_ _05235_ _05238_ _05239_ _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11339_ _00381_ _01524_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12107__A4 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07166__C _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07519__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13009_ _05812_ _05813_ _05912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06880_ _05647_ _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XPHY_EDGE_ROW_145_Left_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08550_ _06642_ _00370_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12815__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07501_ _00505_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08481_ _01263_ _01379_ _01380_ _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_102_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07432_ _05822_ _00446_ _00447_ _00448_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_92_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08247__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07363_ DDS_Stage.LCU.state\[0\] _00400_ DDS_Stage.LCU.SelMuxConfig _00401_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_85_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13240__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09102_ _01916_ _01919_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_154_Left_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09995__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07294_ _05658_ _06232_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_127_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09033_ _01924_ _01925_ _01926_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_115_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12200__B1 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11554__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09935_ _02808_ _02818_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11306__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09866_ _02644_ _02652_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08817_ _06659_ _00370_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09797_ _02647_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_146_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07930__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08748_ _01564_ _01643_ _01644_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08679_ _06308_ _00398_ _00394_ net152 _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_68_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10710_ _03567_ _03583_ _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_49_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11690_ _04531_ _04532_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_83_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10641_ _03435_ _03439_ _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09435__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13360_ _06204_ _06208_ _06291_ _06292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10572_ _03287_ _03375_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07997__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12990__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12311_ _05101_ _05102_ _05155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13291_ _06215_ _06212_ _06216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_121_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12242_ _05037_ _05046_ _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06950__I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12173_ _04944_ _05015_ _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_82_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11124_ _03950_ _03952_ _03966_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_11055_ _03870_ _03878_ _03897_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10006_ _02880_ _02888_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07921__A1 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11957_ _04799_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_86_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10908_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-17\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-17\]
+ _05171_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11888_ _04538_ _04598_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_55_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13627_ _06577_ _06551_ _06527_ _06578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10839_ _03639_ _03710_ _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13558_ _06462_ _06504_ _06505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11784__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12509_ _03930_ _03946_ _05370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_113_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13489_ _06409_ _06430_ _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_113_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06860__I _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11536__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07177__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08401__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07981_ _00394_ _05833_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06963__A2 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ net96 _06674_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06932_ _05409_ _06211_ _06221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_129_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11839__A3 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09901__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ _02443_ _02537_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06863_ _05442_ _05463_ _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__07912__A1 _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08602_ _01484_ _01486_ _01500_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_96_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09582_ _02370_ _02384_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08533_ _01425_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11472__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08464_ _01274_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_147_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07140__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07415_ _05658_ _00433_ _00434_ _06732_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_46_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08395_ _01293_ _01294_ _01295_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_135_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07346_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-4\] _00388_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XANTENNA__09968__A2 _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12972__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11775__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07277_ _06146_ _00333_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09016_ _01901_ _01909_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06954__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09918_ _02710_ _02713_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08156__A1 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09849_ _02729_ _02733_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_137_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07903__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12860_ _05748_ _05749_ _05750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output35_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11811_ _04653_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12791_ _05662_ _05674_ _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08459__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10266__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11742_ _04570_ _04583_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_96_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11673_ _04466_ _04515_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13412_ _03556_ _00387_ _06347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11215__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10624_ net63 _06738_ net57 _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06890__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13343_ _06272_ _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10555_ _03037_ _03430_ _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08092__B1 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13274_ _06134_ _06198_ _06199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10486_ _03037_ _03280_ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11518__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12225_ _05063_ _05067_ _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12156_ _04989_ _04997_ _04998_ _04999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_112_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11107_ _03837_ _03841_ _03949_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12087_ _04915_ _04928_ _04929_ _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_88_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11038_ _03866_ _03879_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09895__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10151__B _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09647__A1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12989_ _03485_ _00375_ _05890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09647__B2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11454__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06855__I _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07200_ _05387_ _06809_ _06810_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06881__A1 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08180_ _01080_ _01081_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07131_ _05387_ _06747_ _06750_ _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_99_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07062_ _05822_ _06691_ _06692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10326__B net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12706__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08386__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10193__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ _00840_ _00865_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08138__A1 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09703_ _02567_ _02568_ _02588_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06915_ _05864_ _06028_ _05182_ _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07895_ _00792_ _00796_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09634_ net158 _06710_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10496__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06846_ _05280_ net18 net17 _05291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_69_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09565_ _00379_ _06685_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09638__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08516_ _01399_ _01401_ _01415_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_78_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09496_ _02370_ _02384_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07113__A2 _06732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08447_ _01346_ _01230_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_65_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08378_ net143 _06637_ _06633_ net91 _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12945__A1 _05740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07329_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-8\] _00375_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_33_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09810__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10340_ _03124_ _03127_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07529__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _03142_ _03150_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12010_ _04852_ _04848_ _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_100_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10184__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08129__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11279__A4 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12912_ _05710_ _05711_ _05807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07888__B1 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11684__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13892_ _00223_ net36 clknet_leaf_17_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_69_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12843_ _05822_ _05730_ _05731_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_100_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_83_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10239__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11436__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12774_ _05576_ _05589_ _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11725_ _04533_ _04535_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_126_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06863__A1 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11656_ _04472_ _04479_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_154_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10607_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-1\] _03482_ _03414_ _03483_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11587_ _04427_ _04428_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13326_ _06239_ _06253_ _06255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_107_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10538_ _03352_ _03413_ _05182_ _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08080__A3 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13257_ _03340_ _00390_ _06181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10469_ _03257_ _03336_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08368__A1 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12208_ _05050_ _05051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09427__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10175__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13188_ _06050_ _06105_ _06106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06918__A2 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11911__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07040__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12139_ _04882_ _04980_ _04981_ _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13664__A2 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07680_ DDS_Stage.xPoints_Generator1.CosNew\[-4\] _00645_ _00577_ _00646_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ _02239_ _02167_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09096__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08301_ _00934_ _01201_ _01202_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11978__A2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09281_ _02098_ _02127_ _02171_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08232_ _01099_ _01100_ _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ _01047_ _01064_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_132_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07114_ _05658_ _06736_ _06737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10402__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ _00993_ _00994_ _00995_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07045_ _06232_ _05702_ _06555_ _06676_ _06677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__10953__A3 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09020__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06909__A2 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11902__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07031__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08996_ _01834_ _01859_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09308__B1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ net142 _06627_ _06618_ net92 _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_98_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07878_ _00367_ _06523_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08531__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09617_ _02471_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13895__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11418__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09548_ _02431_ _02435_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_65_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07098__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ _02294_ _02297_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08834__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11510_ _04270_ _04283_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_108_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12490_ _05282_ _05350_ _05351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_156_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _04270_ _04283_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11372_ _00384_ _01524_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07259__C _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13111_ _05823_ _05828_ _06023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10323_ _02608_ _02704_ _03201_ _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07270__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13042_ _05867_ _05896_ _05947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10254_ _03060_ _03068_ _03133_ _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09011__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07022__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10185_ _00385_ _06710_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08770__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13646__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13944_ _00275_ net101 clknet_leaf_28_clk net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_89_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13886__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13875_ _00206_ net36 clknet_leaf_55_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_0_88_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12826_ _05708_ _05712_ _05714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07089__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12757_ _05632_ _05637_ _05639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_45_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11708_ _04522_ _04550_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_154_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12688_ _05473_ _05562_ _05563_ _05564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12909__A1 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11639_ _04472_ _04479_ _04481_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08589__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09250__A2 _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13309_ _06154_ _06169_ _06235_ _06236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__13810__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13334__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07013__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08850_ _00394_ _06598_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11896__A1 _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07801_ _00716_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08761__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10163__A4 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08781_ _01673_ _01677_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07732_ net6 DDS_Stage.xPoints_Generator1.RegF\[-2\] _00667_ _00681_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_140_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13877__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07663_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-7\] DDS_Stage.xPoints_Generator1.RegFrequency\[-7\]
+ _00626_ _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10320__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09402_ _06649_ net95 _06710_ net58 _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_88_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07594_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[29\] _00573_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09333_ _02161_ _02163_ _02223_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_TAPCELL_ROW_36_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11415__A4 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09264_ _02134_ _02136_ _02133_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_30_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08215_ _01115_ _01116_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_146_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08029__B1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09195_ _02083_ _02086_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08146_ _01028_ _01032_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13801__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07252__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08077_ _00976_ _00977_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07252__B2 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07028_ _06146_ _06662_ _06663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07004__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08979_ _05387_ _01871_ _01873_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold55 FreqPhase[8] net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold66 net11 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold77 _05346_ net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold88 FreqPhase[14] net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_11990_ _04817_ _04818_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08504__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08504__B2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13868__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10941_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-1\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-1\]
+ _05171_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10311__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13660_ _05442_ _05387_ _00568_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10872_ _03647_ _03709_ _03742_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12611_ _03485_ net148 _00361_ _00365_ _05480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_155_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13591_ _06493_ _06494_ _06540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12603__A3 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12542_ _05374_ _05391_ _05404_ _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_136_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07491__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12473_ _05235_ _05238_ _05328_ _05331_ _05239_ _05332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_81_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07618__I0 DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_11424_ _00361_ _02153_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07243__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11355_ _04196_ _04197_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_132_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12119__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08991__A1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10306_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-5\] _03185_ _03186_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11286_ _00361_ _02854_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13025_ _05823_ _05828_ _05929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10237_ _03115_ _03116_ _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11878__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08743__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10168_ _03030_ _03048_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_109_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _02904_ _02905_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13859__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13927_ _00258_ net36 clknet_leaf_29_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_77_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13858_ _00189_ net36 clknet_leaf_49_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_92_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12809_ _05602_ _05611_ _05694_ _05695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13789_ _00120_ net36 clknet_leaf_63_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_18_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09471__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10081__A3 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08000_ _00900_ _00901_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_100_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_5__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07234__A1 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09951_ _02687_ _02747_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08902_ _01770_ _01773_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_111_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09882_ _02744_ _02745_ _02765_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08833_ _01646_ _01727_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08764_ _00394_ net156 _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07715_ _00672_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_49_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11097__A2 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08695_ net60 _06659_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07646_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-9\] _00616_ _00395_ _00617_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_146_Right_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12046__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07577_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[22\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-9\]
+ _00395_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09316_ _02119_ _02205_ _02206_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09462__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_153_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09247_ _02055_ _02062_ _02138_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__07473__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _01994_ _02012_ _02069_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_32_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09214__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08129_ net73 _06416_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07225__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput23 net23 Cos_Out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11140_ _03930_ _03946_ _03982_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput34 net34 Cos_Out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_73_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11071_ _03882_ _03912_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10022_ _00385_ _06701_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12521__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11973_ _00369_ _02584_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10135__I1 _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13712_ _00047_ clknet_leaf_13_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10924_ _03778_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10835__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13643_ _06536_ _06537_ _06595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10855_ _05822_ _03724_ _03726_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13574_ _06470_ _06503_ _06521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10786_ _03654_ _03658_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_30_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_9_clk_I clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08256__A3 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07464__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12525_ _03340_ _00365_ _05386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12456_ _03763_ _05310_ _05314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11407_ _04245_ _04249_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11012__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12387_ _04872_ _04942_ _05239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_23_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11338_ _00384_ _01430_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10771__A1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10154__B _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07447__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11269_ _00381_ _00384_ _02409_ _02238_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_120_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07519__A2 _06623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13008_ _05812_ _05813_ _05911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11720__B1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07463__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07500_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-7\] _00502_ _00504_
+ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09141__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08480_ _01264_ _01265_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07431_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-19\] _00448_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07362_ DDS_Stage.LCU.state\[2\] _05226_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09101_ _01901_ _01909_ _01993_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_116_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07455__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07293_ _05409_ _06555_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09032_ net95 _06633_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07207__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12200__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12200__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08955__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09934_ _02811_ _02817_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09865_ _02644_ _02652_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11711__B1 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08816_ _01708_ _01711_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09796_ _02673_ _02675_ _02680_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_0_84_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07930__A2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13706__CLK clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08747_ _01565_ _01566_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08678_ _01496_ _01498_ _01575_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07629_ _00600_ _00601_ _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10640_ _03311_ _03456_ _03514_ _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09435__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07446__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10571_ _03371_ _03374_ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07446__B2 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12310_ _05150_ _05151_ _05153_ _05154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_51_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07997__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12990__A2 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13290_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-5\] _06209_ _06215_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_23_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09199__A1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12241_ _05083_ _05071_ _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_75_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12172_ _04985_ _05013_ _05014_ _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11123_ _03960_ _03965_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11054_ _03873_ _03877_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10005_ _02792_ _02887_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09371__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07921__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11956_ _04794_ _04798_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_86_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10907_ _05387_ _03768_ _03769_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11887_ _04644_ _04698_ _04729_ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_129_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13626_ _06528_ _06577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10838_ _03647_ _03709_ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07437__A1 _06698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10769_ _02704_ _03640_ _03641_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_13557_ _06470_ _06503_ _06504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07437__B2 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11784__A3 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12508_ _05365_ _05368_ _05369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13488_ _06411_ _06429_ _06430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_117_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12439_ _04740_ _04741_ _05209_ _05294_ _05295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_124_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07980_ _00858_ _00881_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06931_ _05420_ _05442_ _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__11839__A4 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09650_ _02533_ _02536_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06862_ _05452_ _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_59_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08601_ _01494_ _01499_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07912__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09581_ _02419_ _02468_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09114__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08532_ _01427_ _01429_ _01431_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08463_ _01361_ _01362_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11472__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07414_ _05658_ _06705_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08394_ _05864_ _00394_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07428__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07345_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-4\] _00387_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_18_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_clk clknet_3_5__leaf_clk clknet_leaf_30_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12972__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07276_ _05995_ _06622_ _00332_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09015_ _01904_ _01908_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_130_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09917_ _02726_ _02734_ _02800_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08156__A2 _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09848_ _02730_ _02731_ _02732_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__07903__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09779_ _02494_ _02661_ _02664_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09105__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11810_ _04652_ _04650_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12790_ _05668_ _05673_ _05674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07323__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11741_ _04570_ _04583_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11672_ _04513_ _04514_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10623_ _03432_ _03441_ _03497_ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13411_ _06345_ _06346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07419__A1 _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11215__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07419__B2 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06890__A2 _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_21_clk clknet_3_7__leaf_clk clknet_leaf_21_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13342_ _06187_ _06270_ _06271_ _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10554_ net57 _02704_ _03429_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08092__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08092__B2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13273_ _06197_ _06198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10485_ _03282_ _03290_ _03361_ _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12224_ _05066_ _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10726__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12155_ _04993_ _04996_ _04998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_112_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11106_ _03842_ _03844_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12086_ _04926_ _04927_ _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09344__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11037_ _03866_ _03879_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_88_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11151__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09895__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12988_ net147 _00378_ _05889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09647__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11454__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11939_ _04781_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13609_ _06557_ _06558_ _06559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06881__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_12_clk clknet_3_3__leaf_clk clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07130_ _05431_ _06566_ _06749_ _06146_ _06750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_131_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08083__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10965__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07061_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-4\] _06691_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07830__A1 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12706__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08386__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10193__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07963_ _00842_ _00864_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_52_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08138__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06914_ _05658_ _05962_ _06017_ _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09702_ _02587_ _02566_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07894_ _00793_ _00794_ _00795_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09633_ _00357_ _06730_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06845_ _05269_ _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XANTENNA__10496__A3 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clone57_I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09564_ _00373_ _06696_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09638__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08515_ _01406_ _01414_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_26_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09495_ _02375_ _02383_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_33_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08446_ _01338_ _01341_ _01344_ _01345_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA_clkbuf_leaf_34_clk_I clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08377_ _00898_ _00903_ _01277_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_92_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07328_ _00374_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09810__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_49_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07821__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ _06491_ _00317_ _00318_ _06629_ _05171_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_60_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10270_ _03145_ _03149_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09023__B1 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09574__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10184__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08129__A2 _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12911_ _05802_ _05805_ _05806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07888__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12881__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07888__B2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11684__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13891_ _00222_ net36 clknet_leaf_11_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_12842_ _05280_ net30 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_83_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11436__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12773_ _05560_ _05575_ _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11724_ _04553_ _04566_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07360__I0 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11655_ _04496_ _04497_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06863__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10606_ _03410_ _03412_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11586_ _04427_ _04428_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10947__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13325_ _06241_ _06252_ _06253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10537_ _03352_ _03413_ _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_114_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08080__A4 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10468_ _02849_ _02930_ _03096_ _03098_ _03099_ _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_13256_ _03266_ _00393_ _06180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08368__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09565__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12207_ _05021_ _05023_ _05049_ _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13187_ _06052_ _06104_ _06105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10399_ _03037_ _03202_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_94_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11372__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10175__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12138_ _04883_ _04884_ _04981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09317__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12069_ _04907_ _04911_ _04912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_1_clk clknet_3_2__leaf_clk clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07879__A1 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12624__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08300_ _00935_ _00936_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11978__A3 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09280_ _02101_ _02126_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07351__I0 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08231_ _01124_ _01132_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_144_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13917__CLK clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08056__A1 _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08162_ _01024_ _01063_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07113_ _05409_ _06732_ _06735_ _06736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11060__B1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08093_ net61 net60 _05833_ _05398_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07803__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07044_ _05518_ _06340_ _06676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10953__A4 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11902__A3 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08995_ _01887_ _01888_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09308__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09308__B2 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07946_ _00811_ _00816_ _00847_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11115__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ _00357_ _06618_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_98_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08531__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09616_ _02414_ _02478_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11418__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09547_ _02432_ _02433_ _02434_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_65_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09478_ _02263_ _02271_ _02366_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_109_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08429_ _01069_ _01094_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08047__A1 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11440_ _04273_ _04282_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11371_ _04183_ _04212_ _04213_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10322_ net63 _06710_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13110_ _05829_ _05928_ _06022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_132_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13041_ _05942_ _05945_ _05946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10253_ _03063_ _03132_ _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10157__A2 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11354__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10184_ _00388_ _06708_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08770__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13943_ _00274_ net101 clknet_leaf_29_clk net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_88_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13874_ _00205_ net36 clknet_leaf_60_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_69_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12606__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12825_ _05709_ _05710_ _05711_ _05712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_57_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12756_ _05632_ _05637_ _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11707_ _04521_ _04523_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12687_ net87 _00354_ _03558_ _03679_ _05563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_37_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12909__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11638_ _04477_ _04480_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13031__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08589__A2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11569_ _04345_ _04411_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_80_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11593__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13308_ _06150_ _06153_ _06235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13334__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13239_ _06159_ _06160_ _06161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_126_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11345__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07800_ _00355_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[17\] _00395_ _00716_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08761__A2 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08780_ _01674_ _01675_ _01676_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07731_ _00680_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_140_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07662_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-7\] DDS_Stage.xPoints_Generator1.RegFrequency\[-7\]
+ _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_140_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09401_ _02277_ _02290_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07593_ _05387_ _00571_ _00572_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_105_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09332_ _02170_ _02222_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10084__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11281__B1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09263_ _06059_ _02152_ _02154_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_146_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08214_ _00988_ _01036_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08029__A1 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08029__B2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09194_ _02084_ _02085_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_138_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08145_ _01044_ _01045_ _01046_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11584__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08076_ _00976_ _00977_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_114_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07027_ _05583_ _06211_ _06661_ _06662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_11_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08201__A1 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07004__A2 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08978_ _01872_ _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold56 net15 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold67 net121 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold78 _00290_ net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07929_ _06308_ _00382_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold89 FreqPhase[12] net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08504__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10940_ _03786_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07563__I0 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10871_ _03642_ _03708_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12610_ _03340_ _00369_ _05479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13590_ _06538_ _06539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12603__A4 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12541_ _05394_ _05403_ _05404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13013__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12472_ _05329_ _05288_ _05330_ _05331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07491__A2 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11423_ _00365_ _02051_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11575__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11354_ _00361_ _01956_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10305_ _03090_ _03093_ _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08991__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11285_ _00369_ _02586_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_91_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10236_ _03034_ _03037_ _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_5_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_91_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13024_ _05926_ _05927_ _05928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11878__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10925__I1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08743__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _03039_ _03047_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_109_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10098_ _02976_ _02979_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13926_ _00257_ net36 clknet_leaf_28_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_92_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13857_ _00188_ net36 clknet_leaf_51_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_53_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12808_ _05606_ _05693_ _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13788_ _00119_ net36 clknet_leaf_63_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12739_ _05455_ _05527_ _05620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13004__A1 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13795__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07196__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09950_ _02766_ _02833_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06993__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-19\] _01796_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09881_ _02764_ _02743_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08832_ _01647_ _01648_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08763_ _00398_ net153 _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07714_ net118 DDS_Stage.xPoints_Generator1.RegF\[-11\] _00667_ _00672_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_49_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08694_ net91 _06654_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13661__B _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07645_ DDS_Stage.xPoints_Generator1.CosNew\[-9\] _00615_ _00577_ _00616_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07576_ _00562_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12046__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09998__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09315_ net61 net60 _06685_ _06691_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_118_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09246_ _02133_ _02137_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_118_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09177_ _01997_ _02011_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_90_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ net158 _06179_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07225__A2 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13786__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08059_ _00957_ _00960_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xoutput24 net24 Cos_Out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 net35 Cos_Out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06984__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11070_ _03882_ _03912_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_73_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10021_ _00388_ _06696_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09922__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07553__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13482__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11972_ _04804_ _04813_ _04814_ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13711_ _00046_ clknet_3_5__leaf_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10923_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-10\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-10\]
+ _05171_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13642_ _06532_ _06592_ _06593_ _06594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10854_ _05280_ _03725_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13573_ _06472_ _06501_ _06520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10785_ _03592_ _03657_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_30_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08256__A4 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12524_ _03266_ _00369_ _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07464__A2 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12455_ _03763_ _05310_ _05311_ _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_34_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06913__B _06006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11406_ _04246_ _04247_ _04248_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_62_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12386_ _05014_ _05236_ _04944_ _05238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_50_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11337_ _04179_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10771__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11268_ _04110_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08177__B1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13007_ _05905_ _05909_ _05910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10219_ _02758_ _02850_ _03096_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_11199_ _04039_ _04040_ _04041_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11720__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11720__B2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13473__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09141__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13909_ _00240_ net36 clknet_leaf_24_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[31\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_18_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07152__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07430_ _06232_ _06756_ _06820_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11236__B1 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07361_ _00399_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11787__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09100_ _01904_ _01908_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07292_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[1\] _00346_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_128_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09031_ net138 _06696_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_135_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07207__A2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12200__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08955__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06966__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09933_ _02815_ _02816_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09904__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09864_ _02684_ _02748_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11711__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11711__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08815_ _01709_ _01710_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10080__B _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09795_ _02576_ _02577_ _02676_ _02678_ _02679_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13940__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07930__A3 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08746_ _01565_ _01566_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_77_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07143__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08677_ net137 net96 net152 _06672_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_68_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07628_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-12\] DDS_Stage.xPoints_Generator1.RegFrequency\[-12\]
+ _00596_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07559_ _00350_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_153_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10570_ _03311_ _03392_ _03445_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_146_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07446__A2 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09229_ net60 _06691_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12240_ _05078_ _05082_ _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09199__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12171_ _05011_ _05012_ _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06957__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11122_ _03961_ _03964_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11053_ _03885_ _03895_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_101_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11702__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10004_ _02883_ _02886_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09371__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13931__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11955_ _04797_ _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07134__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10906_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-18\] _03769_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08882__A1 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13207__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11886_ _04614_ _04643_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13625_ _06524_ _06561_ _06574_ _06575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10837_ _03642_ _03708_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_13_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13556_ _06472_ _06501_ _06503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10768_ net58 net63 _06744_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_55_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12507_ _04019_ _04020_ _05367_ _05368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13487_ _06418_ _06428_ _06429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11784__A4 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10699_ _03571_ _03572_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12438_ _05242_ _05243_ _05294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12369_ _05217_ _05218_ _05219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06930_ _06059_ _06168_ _06190_ _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06861_ DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[1\] _05452_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__13922__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08600_ _01497_ _01498_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09580_ _02446_ _02467_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09114__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08531_ _05280_ _01430_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07125__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08462_ _06637_ _00370_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07413_ _05507_ _06788_ _00341_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10680__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08393_ _00398_ _05833_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07344_ _00386_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07275_ _06232_ _06645_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09014_ _01905_ _01906_ _01907_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_103_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12185__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13386__B _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09916_ _02729_ _02733_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_8_clk_I clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ _00385_ _06691_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13913__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07903__A3 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09778_ _02663_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09105__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08729_ _06642_ _00373_ _01559_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_1_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07116__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11740_ _04574_ _04582_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_68_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11671_ _04464_ _04465_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13410_ _06274_ _06343_ _06344_ _06345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10622_ _03428_ _03431_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13341_ _06188_ _06189_ _06271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10553_ net63 _06738_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08092__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13272_ _06143_ _06196_ _06197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10484_ _03278_ _03281_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12223_ _05056_ _05064_ _05065_ _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11923__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12154_ _04993_ _04996_ _04997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_112_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11105_ _03918_ _03947_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12085_ _04926_ _04927_ _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11036_ _03870_ _03878_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_88_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13904__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11151__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07514__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12987_ _05771_ _05885_ _05887_ _05888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07107__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12100__A1 _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11938_ _04748_ _04750_ _04780_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08855__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11869_ _04707_ _04711_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13608_ _03485_ _00397_ _06487_ _06558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_55_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13539_ _03485_ _00397_ _06484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08083__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10965__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07060_ _05658_ _06689_ _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07830__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09032__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07962_ _00846_ _00863_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_52_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09701_ _02564_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06913_ _05409_ _05984_ _06006_ _05658_ _06017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07893_ net143 _06618_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09632_ _02427_ _02517_ _02518_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06844_ _05171_ _05269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10496__A4 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09563_ _02449_ _02450_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08514_ _01409_ _01413_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09494_ _02378_ _02382_ _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_33_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ _01218_ _01223_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08376_ _00893_ _00897_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10405__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ _00372_ _00373_ _05182_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09810__A3 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07258_ _06146_ _06623_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07189_ _06801_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09023__A1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09023__B2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11905__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09574__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13658__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07188__I1 _06800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12910_ _05803_ _05804_ _05805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07888__A2 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13890_ _00221_ net36 clknet_leaf_36_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__12881__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12841_ _05727_ _05729_ _05730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12772_ _05591_ _05613_ _05653_ _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10644__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11723_ _04560_ _04565_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07360__I1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11654_ _04442_ _04450_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10605_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[0\] _03472_ _03480_ _03481_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_37_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07289__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09262__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11585_ _00361_ _01794_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10947__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13324_ _06244_ _06251_ _06252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_hold65_I FreqPhase[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10536_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-1\] _03410_ _03412_ _03413_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_114_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12149__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13255_ _03189_ _00397_ _06178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10467_ _02681_ _03343_ _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06921__B _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12206_ _00381_ _00384_ _01794_ _01792_ _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_86_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09565__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13186_ _06079_ _06102_ _06104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10398_ _03204_ _03212_ _03275_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_94_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11372__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12137_ _04883_ _04884_ _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12068_ _04910_ _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11019_ _03859_ _03860_ _03861_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_95_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07879__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_125_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08828__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12624__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10635__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11978__A4 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07500__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07351__I1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08230_ _01125_ _01131_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _01062_ _01049_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08056__A2 _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07112_ _05409_ _06734_ _06735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11060__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08092_ net60 _05833_ _05398_ net61 _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07803__A2 _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11060__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07043_ _06059_ _06640_ _06675_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09005__A1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11902__A4 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08994_ _00370_ _06672_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09308__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07945_ _00806_ _00810_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13664__B _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11115__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone9_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07876_ _00775_ _00776_ _00777_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09615_ _02416_ _02477_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10874__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09546_ net137 _06738_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10626__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09477_ _02266_ _02270_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09492__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08428_ _01315_ _01322_ _01324_ _01325_ _01327_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_19_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08047__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08359_ _00914_ _00915_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_117_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07255__B1 _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11370_ _04181_ _04182_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_62_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10321_ _03115_ _03199_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13040_ _05943_ _05944_ _05945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10252_ _03067_ _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11354__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10183_ _00382_ _06724_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08507__B1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13942_ _00273_ net101 clknet_leaf_29_clk net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13873_ _00204_ net36 clknet_leaf_64_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_12824_ _03189_ _00381_ _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12606__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12755_ _05360_ _05633_ _05636_ _05637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09483__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11706_ _04544_ _04548_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_126_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12686_ _00354_ _03558_ _03679_ net87 _05562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_127_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11637_ _04478_ _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_86_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08589__A3 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11568_ _04352_ _04410_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_96_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11593__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13307_ _06171_ _06194_ _06233_ _06234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10519_ _03360_ _03395_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11499_ _04321_ _04341_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13238_ _00369_ _03725_ _06060_ _06160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07466__C _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07549__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11345__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13169_ _05965_ _05975_ _06085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_clk_I clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08761__A3 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07730_ net5 DDS_Stage.xPoints_Generator1.RegF\[-3\] _00667_ _00680_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07661_ _00629_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_140_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_48_clk_I clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09400_ _02285_ _02289_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07592_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-3\] _05182_ _00572_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07702__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09331_ _02172_ _02221_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11805__B1 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_47_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10084__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11281__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09262_ _05280_ _02153_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11281__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08213_ _01098_ _01113_ _01114_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08029__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09193_ _00376_ _06672_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11033__A1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08144_ _01020_ _01034_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12781__A1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11584__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08075_ _00769_ _00867_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_151_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07026_ _05409_ _05420_ _05474_ _06661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_140_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08201__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08977_ _01868_ _01870_ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xhold57 FreqPhase[10] net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07928_ _00829_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold68 net10 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold79 net165 net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_39_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07859_ _00757_ _00759_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10870_ _03739_ _03740_ _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09529_ _02356_ _02364_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12540_ _05397_ _05402_ _05403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_109_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12471_ _05211_ _05221_ _05330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13013__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11422_ _00369_ _01956_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11024__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11575__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11353_ _00365_ _01794_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10304_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-4\] _03183_ _03184_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_120_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11284_ _04122_ _04126_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12524__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13023_ _05850_ _05851_ _05925_ _05927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_10235_ net61 net60 net161 _06744_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__11878__A3 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10166_ _02966_ _03046_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_109_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10097_ _02977_ _02978_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13925_ _00256_ net36 clknet_leaf_33_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_107_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13856_ _00187_ net36 clknet_leaf_51_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_122_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12807_ _05610_ _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13787_ DDS_Stage.LCU.SelMuxConfig net36 clknet_leaf_72_clk DDS_Stage.LCU.SelMuxConfigReg
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10999_ _03837_ _03841_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_85_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12738_ _05544_ _05618_ _05619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XPHY_EDGE_ROW_106_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12669_ _05822_ net29 _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13004__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08900_ _05822_ _01794_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06993__A2 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09880_ _02741_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08195__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08831_ _01647_ _01648_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_100_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08762_ _01584_ _01657_ _01658_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07713_ _00671_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08693_ net73 _06664_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07644_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-9\] DDS_Stage.xPoints_Generator1.RegFrequency\[-9\]
+ _00614_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_124_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07575_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[21\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-10\]
+ _00395_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_62_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ net61 _06685_ _06691_ net60 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09998__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09245_ _02134_ _02136_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09176_ _02066_ _02067_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ _00363_ _06308_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07225__A3 _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_133_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08058_ _00958_ _00959_ _00775_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
Xoutput25 net25 Cos_Out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12506__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07009_ _05409_ _06644_ _06646_ _06647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_73_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10020_ _00382_ _06708_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09922__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11971_ _04808_ _04812_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13482__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13710_ _00045_ clknet_leaf_33_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11493__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10922_ _03777_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13641_ _06533_ _06550_ _06593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10853_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[30\] _03725_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_128_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13572_ _06517_ _06518_ _06519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10784_ _03655_ _03656_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08110__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12523_ _05379_ _05383_ _05384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_54_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__A3 _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12454_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-23\] _05296_ _05311_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11405_ _00361_ _02051_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06913__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12385_ _04984_ _05210_ _05236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11336_ _04176_ _04177_ _04178_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11267_ _04107_ _04108_ _04109_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08177__A1 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13006_ _05906_ _05907_ _05909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08177__B2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10218_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-6\] _03097_ _03099_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_11198_ _00381_ _00384_ _02409_ _02238_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__11720__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10149_ _03028_ _03029_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13473__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13908_ _00239_ net36 clknet_leaf_24_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_18_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13839_ _00170_ clknet_leaf_68_clk DDS_Stage.xPoints_Generator1.RegP\[-9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11236__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07360_ _00397_ _00398_ _00395_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11236__B2 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11787__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07291_ _00344_ _00345_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09030_ _00355_ _06691_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_135_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09601__A1 _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08955__A3 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06966__A2 _06576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09932_ _02813_ _02814_ _02812_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09904__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09863_ _02687_ _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_55_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11711__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08814_ _06649_ _00373_ _01641_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_99_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09794_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-10\] _02677_ _02679_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08745_ _01638_ _01641_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_146_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07930__A4 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09668__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08676_ _01484_ _01572_ _01573_ _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07143__A2 _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07627_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-12\] DDS_Stage.xPoints_Generator1.RegFrequency\[-12\]
+ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07558_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[4\] _00552_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_49_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12975__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07489_ _06232_ _06070_ _00455_ _05658_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_63_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09228_ net91 _06685_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12727__A1 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09159_ _05280_ _02051_ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_75_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12170_ _05011_ _05012_ _05013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10202__A2 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11121_ _03962_ _03963_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11052_ _03888_ _03894_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07906__A1 _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10003_ _02884_ _02885_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11702__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09659__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11954_ _04787_ _04795_ _04796_ _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07134__A2 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10905_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-18\] _03768_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_86_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11885_ _04703_ _04719_ _04726_ _04727_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__08882__A2 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13624_ _06467_ _06562_ _06574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10836_ _00398_ _03646_ _03707_ _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07800__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13555_ _06478_ _06500_ _06501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10767_ net58 net63 _06744_ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_43_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12506_ _00397_ _02409_ _04021_ _05367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_13486_ _06422_ _06426_ _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_23_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10698_ _00398_ _00394_ _06738_ _06742_ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_23_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12437_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-20\] _05290_ _05292_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-21\]
+ _05293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_152_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13391__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12368_ _04986_ _05009_ _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07070__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11319_ _04147_ _04160_ _04161_ _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12299_ _05027_ _05141_ _05142_ _05143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06860_ _05431_ _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_98_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08570__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08530_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[2\] _01430_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07490__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07125__A2 _06668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08461_ _01357_ _01360_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07412_ _05387_ _00428_ _00432_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11209__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06884__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08392_ _00900_ _01292_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__07710__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07343_ _00384_ _00385_ _05182_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07274_ _06651_ _00330_ _06759_ _05431_ _06146_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_61_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ _06642_ _00385_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12185__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09915_ _02797_ _02798_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_148_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11696__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09846_ _00388_ _06685_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08561__A1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07903__A4 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09777_ _02484_ _02662_ _02573_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06989_ _05583_ _06469_ _06630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13437__A2 _06374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08728_ _01557_ _01558_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_1_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07116__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08659_ _06633_ _00379_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06875__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11670_ _04507_ _04511_ _04512_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_138_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10621_ _03443_ _03458_ _03495_ _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09813__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13340_ _06188_ _06189_ _06270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10552_ _03115_ _03427_ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13271_ _06145_ _06195_ _06196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_107_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10483_ _03292_ _03313_ _03359_ _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12222_ _05057_ _05058_ _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_106_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11384__B1 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11923__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07052__A1 _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12153_ _04994_ _04995_ _04917_ _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_102_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11104_ _03930_ _03946_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12084_ _04804_ _04813_ _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11035_ _03877_ _03873_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_88_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12986_ _05772_ _05773_ _05887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_99_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07107__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12100__A2 _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11937_ _00381_ _00384_ _02236_ _02153_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08855__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06866__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11868_ _04708_ _04709_ _04710_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10819_ _03592_ _03657_ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13607_ _06485_ _06486_ _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_55_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11799_ _04639_ _04640_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13538_ _06482_ _06403_ _06483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_99_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07291__A1 _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13469_ _06346_ _06350_ _06408_ _06409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13364__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09032__A2 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07043__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13116__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07961_ _00848_ _00862_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09700_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[16\] _02586_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_52_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06912_ _05420_ _05886_ _05995_ _05409_ _06006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__11678__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07892_ net158 _06598_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09631_ net91 net142 _06708_ _06710_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06843_ DDS_Stage.LCU.state\[1\] _05160_ net125 _05248_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_136_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09562_ _02296_ _02363_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08513_ _01410_ _01411_ _01412_ _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_136_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09493_ _02379_ _02380_ _02381_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10102__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08444_ _01234_ _01342_ _01343_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08375_ _00888_ _00905_ _01275_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10405__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07326_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-9\] _00373_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_16
XANTENNA__11602__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07282__A1 _06081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09810__A4 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07257_ _05658_ _00316_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07188_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-18\] _06800_ _05182_ _06801_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09023__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11366__B1 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11905__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07034__A1 _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13658__A2 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13898__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09829_ _02710_ _02713_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12840_ _05728_ _05639_ _05729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12771_ _05652_ _05590_ _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06848__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11722_ _04561_ _04564_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10644__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11841__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11653_ _04492_ _04494_ _04495_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10604_ _03476_ _03479_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_153_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11584_ _00365_ _01792_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09262__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13323_ _06249_ _06250_ _06251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_80_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07273__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10535_ _03328_ net69 _03411_ _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_114_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12149__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13346__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13254_ _06175_ _06074_ _06176_ _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10466_ _03342_ _03100_ _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_32_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12205_ _05037_ _05046_ _05047_ _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07025__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13185_ _06083_ _06086_ _06101_ _06102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_20_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10397_ _03200_ _03203_ _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_94_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12136_ _04959_ _04977_ _04978_ _04979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12067_ _04754_ _04908_ _04909_ _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11018_ net83 _03189_ _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13889__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12969_ _05770_ _05775_ _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08828__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06839__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08160_ _01061_ _01054_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10399__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ _05908_ _06733_ _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13813__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07264__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08091_ net73 _05864_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11060__A2 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07042_ _05822_ _06674_ _06675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09005__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07016__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11899__A1 _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08764__A1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08993_ _01884_ _01886_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07944_ _00844_ _00845_ _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07875_ net92 net143 _06416_ net156 _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10323__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09614_ _02486_ _02494_ _02484_ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_97_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12076__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09545_ _06664_ net96 _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09476_ _02340_ _02356_ _02364_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_148_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09492__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08427_ _01326_ _01313_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_156_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08358_ _00858_ _00881_ _00885_ _00886_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_156_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13804__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07255__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07309_ _05280_ net70 _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08289_ _01181_ _01190_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_117_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10320_ _03037_ _03119_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07007__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10251_ _03114_ _03130_ _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10182_ _02984_ _03061_ _03062_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08507__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13500__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08507__B2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13941_ _00272_ net101 clknet_leaf_29_clk net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_13872_ _00203_ net36 clknet_leaf_50_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_12823_ _03018_ _00384_ _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11814__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12754_ _05634_ _05635_ _05636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09483__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11705_ _04545_ _04546_ _04547_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_12685_ _05478_ _05483_ _05559_ _05560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13567__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11636_ _04477_ _04478_ _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07246__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11567_ _04409_ _04355_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_52_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08589__A4 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08994__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10518_ _03378_ _03394_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13306_ _06149_ _06170_ _06233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11498_ _04324_ _04326_ _04340_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_97_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13237_ _00361_ _00365_ _03727_ _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10449_ _03191_ _03325_ _03326_ _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13168_ _05968_ _06084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10553__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12119_ _00372_ _02236_ _02153_ _00375_ _04962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13099_ _05854_ _06009_ _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08761__A4 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07660_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-7\] _00628_ _00395_ _00629_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07591_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[28\] _00571_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09330_ _02192_ _02220_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_153_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11805__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11805__B2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09261_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[10\] _02153_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07485__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10084__A3 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11281__A2 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08212_ _01111_ _01112_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09192_ _06664_ _00379_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08143_ _01020_ _01034_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07237__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12230__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11033__A2 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12781__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08074_ _00947_ _00973_ _00975_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10792__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_151_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07025_ _06059_ _06658_ _06660_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09785__I0 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08976_ _01868_ _01870_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold58 net3 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07927_ _00743_ _00745_ _00828_ _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold69 FreqPhase[3] net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_39_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07858_ _00757_ _00759_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07789_ _00710_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09528_ _02335_ _02388_ _02415_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07476__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ net142 _06708_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13549__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12470_ _05211_ _05221_ _05329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_81_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11421_ _04259_ _04263_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07228__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11024__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11352_ _00369_ _01792_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_78_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10303_ _03182_ _03170_ _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_105_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11283_ _04123_ _04125_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13022_ _05850_ _05851_ _05925_ _05926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_120_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10234_ _03039_ _03047_ _03113_ _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12524__A2 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11878__A4 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _03042_ _03045_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07951__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10096_ _00376_ _06730_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13924_ _00255_ net36 clknet_leaf_32_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_107_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08900__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13855_ _00186_ net36 clknet_leaf_67_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_92_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_122_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12806_ _05657_ _05690_ _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_128_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13786_ _00291_ net36 clknet_leaf_75_clk DDS_Stage.LCU.state\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10998_ _03838_ _03839_ _03840_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_97_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07467__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12737_ _05546_ _05617_ _05618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_32_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12460__B2 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-20\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12668_ _05822_ _05541_ _05542_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11619_ _04460_ _04461_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_12599_ _05391_ _05404_ _05466_ _05467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07477__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10774__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10526__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08195__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09392__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08830_ _01722_ _01725_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08761_ net58 net95 net155 _06674_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07712_ net10 DDS_Stage.xPoints_Generator1.RegF\[-12\] _00667_ _00671_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08692_ _01490_ _01588_ _01589_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_49_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07643_ _00612_ _00613_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07574_ _00561_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09313_ _02115_ _02123_ _02203_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07458__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_60_clk clknet_3_1__leaf_clk clknet_leaf_60_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09244_ _01979_ _02134_ _02135_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_119_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09175_ _01990_ _02043_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08126_ _01012_ _01026_ _01027_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08958__A1 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10765__A1 _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08057_ _06523_ _00362_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xoutput26 net26 Cos_Out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_141_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07008_ _05409_ _05431_ _06645_ _06646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__12506__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09907__B1 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08959_ net143 _06674_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09135__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11970_ _04808_ _04812_ _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_99_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10921_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-11\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-11\]
+ _05171_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12690__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11493__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13640_ _06533_ _06550_ _06592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10852_ _03721_ _03723_ _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07449__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10783_ _03503_ _03574_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13571_ _06459_ _06505_ _06518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12442__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_51_clk clknet_3_1__leaf_clk clknet_leaf_51_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08110__A2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_clk_I clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12522_ _05380_ _05381_ _05382_ _05383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_136_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12453_ _05164_ _05309_ _05310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11404_ _00365_ _01956_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12384_ _04872_ _04942_ _05235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10756__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_47_clk_I clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11335_ _00381_ _00384_ _01430_ _01249_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07621__A1 DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_11266_ _00381_ _00384_ _02238_ _02236_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08177__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13005_ _03018_ _00390_ _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10217_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-7\] _03014_ _03097_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-6\]
+ _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_11197_ _00381_ _02409_ _02238_ _00384_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_94_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10148_ _02961_ _02969_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10079_ _02952_ _02960_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13907_ _00238_ net36 clknet_leaf_24_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[29\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_18_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13838_ _00169_ clknet_leaf_68_clk DDS_Stage.xPoints_Generator1.RegP\[-10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11236__A2 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13769_ _00104_ clknet_leaf_11_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_leaf_42_clk clknet_3_4__leaf_clk clknet_leaf_42_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07290_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[0\] _00345_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10995__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10907__B _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08955__A4 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07708__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09931_ _02812_ _02813_ _02814_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_110_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09862_ _02746_ _02738_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_55_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08813_ _01639_ _01640_ _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09793_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-11\] _02667_ _02677_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-10\]
+ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_139_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08744_ _01639_ _01640_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_146_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09668__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08675_ _01486_ _01500_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07626_ _00599_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07557_ _00550_ _00551_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_33_clk clknet_3_5__leaf_clk clknet_leaf_33_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12975__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07488_ _06753_ _06789_ _00494_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09227_ net73 _06696_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09158_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[9\] _02051_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__12727__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08109_ _00363_ _06179_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_75_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09089_ _01980_ _01981_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07618__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11120_ _00390_ _02499_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06957__A3 _06081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _03890_ _03893_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11163__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07906__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10002_ _00398_ _00394_ _06679_ _06685_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09659__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11953_ _04788_ _04789_ _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10904_ _03767_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_86_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11884_ _04704_ _04718_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13623_ _06516_ _06564_ _06572_ _06573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10835_ _00398_ _00394_ _06744_ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06893__A2 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_clk clknet_3_6__leaf_clk clknet_leaf_24_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08095__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13554_ _06481_ _06499_ _06500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_hold88_I FreqPhase[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10766_ _03031_ _03637_ _03638_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_137_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12505_ _04015_ _05363_ _05364_ _05365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07842__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10697_ _00398_ _06738_ _06742_ _00394_ _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13485_ _06423_ _06424_ _06425_ _06426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_23_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12436_ _05283_ _05287_ _05292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_117_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13391__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12367_ _05128_ _05214_ _05216_ _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11318_ _04158_ _04159_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_121_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12298_ _05028_ _05029_ _05142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11249_ _03866_ _03879_ _03854_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_38_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08570__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12103__B1 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08460_ _01358_ _01359_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07411_ _05387_ _00431_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08391_ _00899_ _00900_ _00901_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11209__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06884__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_clk clknet_3_6__leaf_clk clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07342_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-5\] _00385_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07273_ _05409_ _05431_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09012_ _06637_ _00388_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09914_ _02773_ _02770_ _02796_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_148_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_70_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09845_ _00382_ _06696_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12893__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11696__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08561__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09776_ _02572_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06988_ _05409_ _05778_ _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_69_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08727_ _01552_ _01570_ _01623_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__12645__A1 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09510__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08658_ _06642_ _00373_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07521__B1 _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-14\] DDS_Stage.xPoints_Generator1.RegFrequency\[-14\]
+ _00579_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06875__A2 _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08589_ _06642_ net61 net60 _06649_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_83_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10408__B1 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10620_ _03426_ _03442_ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10959__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09813__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10551_ _03037_ _03366_ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07824__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10482_ _03276_ _03291_ _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13270_ _06171_ _06194_ _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_20_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12221_ _05057_ _05058_ _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11384__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11384__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12152_ _00354_ _02586_ _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11103_ _03932_ _03945_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_112_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12083_ _04916_ _04924_ _04925_ _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11034_ _03874_ _03875_ _03876_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_88_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12985_ _05772_ _05773_ _05885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11936_ _04765_ _04777_ _04778_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06866__A2 _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11867_ net66 net54 _01430_ _01249_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_13606_ _06481_ _06499_ _06554_ _06556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10818_ _03661_ _03665_ _03689_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_151_Left_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11798_ _04639_ _04640_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13537_ _06244_ _06400_ _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_125_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10749_ _03544_ _03616_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13468_ _06342_ _06352_ _06408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12419_ _05264_ _05267_ _05273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_23_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13399_ _06273_ _06278_ _06332_ _06333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07960_ _00856_ _00861_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_4_clk clknet_3_6__leaf_clk clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06911_ _05420_ _05680_ _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07891_ _00357_ _06627_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11678__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_155_Right_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09630_ net91 _06708_ _06710_ net142 _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06842_ _05182_ net18 net17 _05237_ _05248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_143_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09561_ _02359_ _02362_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08512_ net60 _06649_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09492_ _00385_ _06672_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10102__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08443_ _01199_ _01211_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08374_ _00890_ _00904_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07325_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-9\] _00372_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
XFILLER_0_116_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11602__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07256_ _05431_ _05713_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12582__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07187_ _06797_ _06798_ _06799_ _06780_ _06800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_14_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11366__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11366__B2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07034__A2 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11118__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08534__A2 _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09731__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09828_ _02711_ _02712_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09759_ _02545_ _02559_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_69_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12770_ _05558_ _05652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output26_I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07631__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _04562_ _04563_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_25_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11841__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11652_ _04488_ _04491_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10603_ _03405_ _03409_ _03478_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11583_ _00369_ _01693_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13322_ _00378_ _03679_ _06250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07273__A2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10534_ _03324_ _03327_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12149__A3 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13346__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13253_ _06066_ _06076_ _06176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10465_ _03094_ _03184_ _03257_ _03336_ _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_60_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12204_ _05040_ _05045_ _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13184_ _06091_ _06100_ _06101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10396_ _03214_ _03237_ _03273_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_94_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12135_ _04975_ _04976_ _04978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_102_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07806__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12066_ _04755_ _04756_ _04909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11017_ _00351_ _03266_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12968_ _05865_ _05866_ _05867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10096__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11919_ _00372_ _02409_ _02238_ _00375_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12899_ _05777_ _05792_ _05793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09789__A1 _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07110_ _05420_ _05669_ _06733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_83_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ _00991_ _00989_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07041_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-7\] _06674_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_63_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11348__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11899__A2 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10020__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08764__A2 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08992_ _01819_ _01820_ _01885_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07716__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07943_ _00394_ _05398_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09713__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07874_ net92 net153 _06523_ net143 _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10323__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11520__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _06059_ _02498_ _02500_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09544_ _00355_ _06730_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12076__A2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07327__I0 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09475_ _02296_ _02363_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_148_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08426_ _01310_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_93_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08357_ _00917_ _00922_ _01257_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07308_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-13\] _00359_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_150_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07255__A2 _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08288_ _01185_ _01189_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07239_ _06651_ _06714_ _05409_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_132_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11339__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10250_ _03121_ _03129_ _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_14_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07007__A2 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10181_ _02985_ _02986_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_100_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08507__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13940_ _00271_ net101 clknet_leaf_30_clk net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_13871_ _00202_ net36 clknet_leaf_52_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__13740__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07191__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12822_ _02940_ _00387_ _05709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13264__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09468__B1 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12753_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-12\] _05536_ _05538_ _05635_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11814__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11704_ net70 _01693_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12684_ _05472_ _05477_ _05559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08691__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13567__A2 _06512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11635_ _04421_ _04424_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_53_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11578__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07246__A2 _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11566_ _04388_ _04408_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_24_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13305_ _06229_ _06230_ _06231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10517_ _03381_ _03384_ _03393_ _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08994__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11497_ _04334_ _04339_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_123_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13236_ _06071_ _06155_ _06156_ _06158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10448_ _03194_ _03248_ _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10002__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09943__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13167_ _05990_ _05999_ _06082_ _06083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10379_ _03094_ _03184_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10553__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12118_ _00378_ _02051_ _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13098_ _05924_ _06009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_127_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12049_ _04889_ _04891_ _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_140_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07182__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13731__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07590_ _05387_ _00569_ _00570_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13255__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11805__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09260_ _02145_ _02151_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10084__A4 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ _01111_ _01112_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09191_ _00373_ _06674_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08142_ net58 _00355_ net152 net155 _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_60_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07237__A2 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12230__A2 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13798__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08073_ _00970_ _00974_ _00972_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06996__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07024_ _05822_ _06659_ _06660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_151_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09785__I1 _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08975_ _01869_ _01790_ _01783_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07926_ _05864_ _05833_ _00388_ _00385_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xhold48 net102 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold59 FreqPhase[5] net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_39_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07857_ _00739_ _00758_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07173__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07788_ DDS_Stage.xPoints_Generator1.RegFrequency\[-5\] DDS_Stage.xPoints_Generator1.RegF\[-5\]
+ _00402_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06920__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09527_ _02338_ _02387_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09458_ net158 _06701_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13549__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08409_ _01309_ _01251_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09389_ net61 net142 _06691_ _06696_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_136_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11420_ _04260_ _04261_ _04262_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_152_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07228__A2 _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13789__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ _04189_ _04192_ _04193_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_78_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06987__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11980__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10302_ _03171_ _03089_ _03173_ _03179_ _03181_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_104_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11282_ _04122_ _04124_ _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13021_ _05852_ _05854_ _05924_ _05925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10233_ _03032_ _03038_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_91_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11732__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07356__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10164_ _03043_ _03044_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_109_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10095_ _00379_ _06724_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_6_clk_I clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13923_ _00254_ net36 clknet_leaf_33_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_107_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07164__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08900__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13237__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13854_ _00185_ net36 clknet_leaf_67_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_122_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06911__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12805_ _05675_ _05689_ _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13785_ net130 net36 clknet_leaf_75_clk DDS_Stage.LCU.state\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_57_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10997_ _00384_ net135 _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12736_ _05554_ _05615_ _05617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_85_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12667_ _05280_ net28 _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11618_ _04285_ _04286_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_136_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12598_ _05376_ _05390_ _05466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11549_ _04313_ _04317_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10774__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13219_ _06086_ _06101_ _06139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_0_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09392__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13952__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08760_ net95 net155 _06674_ net137 _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_29_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07711_ _00670_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08691_ net61 net60 _06649_ _06654_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07155__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07642_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-10\] DDS_Stage.xPoints_Generator1.RegFrequency\[-10\]
+ _00608_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06902__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07573_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[20\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-11\]
+ _00395_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_62_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09312_ _02118_ _02122_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09243_ _01980_ _01981_ _02044_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_32_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_38_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09174_ _01992_ _02042_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08125_ net61 net142 _06179_ _05864_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08958__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06969__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11962__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08056_ _00367_ _06416_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07007_ _05420_ _05452_ _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xoutput27 net27 Cos_Out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_102_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09907__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09907__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11714__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13943__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08958_ net158 _06672_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09135__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07909_ _00806_ _00810_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08889_ _01613_ _01606_ _01687_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10920_ _05822_ _06824_ _03776_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12690__A2 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10851_ _03722_ _03677_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13570_ _06462_ _06504_ _06517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08646__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10782_ _03570_ _03573_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12442__A2 _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12521_ net86 _03558_ _05382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12452_ _05190_ _05295_ _05308_ _05309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11403_ _00369_ _01794_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12383_ _05231_ _05232_ _05233_ _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_23_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13596__B _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11334_ _00381_ _01430_ _01249_ _00384_ _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_133_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11265_ _00381_ _02238_ _02236_ _00384_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13004_ _02940_ _00393_ _05906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10216_ _03007_ _03012_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_11196_ _00387_ _02236_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13934__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10147_ _02952_ _02960_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13458__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07814__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10078_ _02954_ _02959_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07137__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13906_ _00237_ net36 clknet_leaf_23_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[28\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_18_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13837_ _00168_ clknet_leaf_68_clk DDS_Stage.xPoints_Generator1.RegP\[-11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13768_ _00103_ clknet_leaf_8_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12719_ _02586_ _00397_ _05598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13699_ _00034_ clknet_leaf_54_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10995__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11944__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09930_ _00388_ _06691_ _06696_ _00385_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09861_ _02744_ _02745_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13925__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ _01634_ _01652_ _01707_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07009__B _06646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09792_ _02659_ _02665_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07724__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08743_ _06642_ _00376_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07128__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08674_ _01486_ _01500_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07625_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-12\] _00598_ _00395_ _00599_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07556_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[3\] _00551_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_46_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11632__B1 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07487_ _05995_ _06221_ _06146_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09226_ _02034_ _02116_ _02117_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09157_ _01967_ _02048_ _05182_ _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08108_ net158 _05864_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_75_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09088_ _01889_ _01940_ _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08039_ _00750_ _00755_ _00753_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_55_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11699__B1 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11050_ _03891_ _03892_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13916__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11163__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10001_ _00398_ _06679_ _06685_ _00394_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07119__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12112__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11952_ _04788_ _04789_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10903_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-19\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-19\]
+ _05171_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10674__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_64_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_86_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11883_ _04717_ _04724_ _04725_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_95_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13622_ _06519_ _06563_ _06572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10834_ _03705_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10426__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13553_ _06483_ _06498_ _06499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10765_ _03031_ _03579_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08095__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12504_ _04017_ _04031_ _05364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13484_ _00381_ _03725_ _06425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07842__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10696_ _02704_ _03568_ _03569_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12179__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12435_ _05222_ _05289_ _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_117_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12366_ _05121_ _05122_ _05216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_73_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11317_ _04158_ _04159_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_130_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12297_ _05028_ _05029_ _05141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_120_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11248_ _04076_ _04089_ _04090_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13907__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11179_ _04018_ _04021_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12103__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12103__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07530__A1 _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07410_ _06146_ _00429_ _00430_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08390_ _01286_ _01290_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__11209__A3 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07341_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-5\] _00384_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
XFILLER_0_155_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11090__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07272_ _00329_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_42_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09011_ _06649_ _00382_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09035__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11917__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09913_ _02773_ _02770_ _02796_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_112_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09844_ _02636_ _02727_ _02728_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_clk_I clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12893__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09775_ _02660_ _02574_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06987_ _06059_ _06626_ _06628_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08726_ _01555_ _01569_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08849__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12645__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08657_ _01553_ _01554_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_46_clk_I clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07521__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07608_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-14\] _05822_ _00584_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08588_ _06642_ net61 net60 _06649_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_83_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10408__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10408__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07539_ _00536_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10959__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10550_ _03368_ _03376_ _03425_ _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_81_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07824__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09209_ _02024_ _02099_ _02100_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_20_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10481_ _03356_ _03357_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12220_ _05034_ _05061_ _05062_ _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_44_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11384__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12151_ _00351_ _02762_ _04994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11102_ _03936_ _03944_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_112_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12082_ _04920_ _04923_ _04925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_9_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11033_ net83 _03266_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10895__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12984_ _05785_ _05882_ _05883_ _05884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11935_ _04771_ _04776_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07512__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11866_ net70 _01247_ _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13605_ _06483_ _06498_ _06554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10817_ _03634_ _03660_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11797_ _04553_ _04566_ _04568_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_144_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13536_ _06422_ _06426_ _06479_ _06481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10748_ _03621_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_153_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13467_ _06395_ _06406_ _06407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_36_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ _03544_ _03552_ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12418_ _05257_ _05271_ _05260_ _05272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13398_ _06269_ _06279_ _06332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12349_ _05195_ _04410_ _05196_ _05197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06910_ _05420_ _05973_ _05984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07890_ _00779_ _00790_ _00791_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_52_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11678__A3 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06841_ DDS_Stage.LCU.state\[2\] DDS_Stage.LCU.state\[0\] _05226_ _05237_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_65_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09560_ _02375_ _02383_ _02447_ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_143_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08511_ _06642_ net91 _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09491_ _06664_ _00388_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07503__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08442_ _01199_ _01211_ _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08373_ _01258_ _01273_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_46_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07324_ _00371_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11063__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11602__A3 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07255_ _05387_ _00312_ _00313_ _00315_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_143_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07186_ _05409_ _06651_ _06340_ _06799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_42_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11366__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11118__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07990__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10877__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09827_ _00398_ _00394_ _06672_ _06674_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09731__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09758_ _02593_ _02643_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08709_ _01605_ _01533_ _01534_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_96_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09689_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-12\] _02495_ _02576_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_83_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11720_ _00361_ _01693_ _01610_ _00365_ _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11651_ _04474_ _04493_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09247__A1 _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10602_ _03411_ _03477_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11582_ _04421_ _04424_ _04422_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13321_ _06247_ _06248_ _06249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10533_ _03405_ _03409_ _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13252_ _06069_ _06175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12149__A4 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10464_ _05822_ _03339_ _03341_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12203_ _05040_ _05045_ _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13183_ _06095_ _06099_ _06100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10395_ _03198_ _03213_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12134_ _04975_ _04976_ _04977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_94_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07981__A1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12065_ _04755_ _04756_ _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11016_ _00359_ _03018_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_125_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12967_ _05777_ _05792_ _05866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06946__B _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11918_ _00378_ _02236_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10096__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12898_ _05781_ _05791_ _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11849_ _04690_ _04691_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12793__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13519_ _06460_ _06461_ _06462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07040_ _06059_ _06671_ _06673_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11348__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10020__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08991_ _06659_ _00373_ _01821_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_10_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07942_ _00813_ _00814_ _00843_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_76_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09713__A2 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07873_ _00357_ _06598_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11520__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ _05280_ _02499_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07732__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09543_ _02426_ _02430_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_149_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12076__A3 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07327__I1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone48_I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09474_ _02359_ _02362_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_65_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08425_ _01241_ _01242_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_65_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09229__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08356_ _00912_ _01256_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07307_ net161 _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_61_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08287_ _01188_ _01187_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_116_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07238_ _05822_ _00298_ _00300_ _00301_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__11339__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12536__A1 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07169_ _05550_ _06681_ _06373_ _05658_ _06784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_131_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10180_ _02985_ _02986_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_100_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13870_ _00201_ net36 clknet_leaf_53_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07191__A2 _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12821_ _05607_ _05706_ _05707_ _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09468__B2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13264__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11275__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12752_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-12\] _05536_ _05634_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11703_ net54 _01792_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12683_ _05486_ _05500_ _05557_ _05558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08691__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11634_ _04473_ _04476_ _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_53_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11578__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11565_ _04391_ _04393_ _04407_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09640__A1 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_96_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold63_I FreqPhase[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13304_ _06224_ _06225_ _06228_ _06230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_10516_ _03311_ _03392_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_134_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11496_ _04335_ _04338_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13235_ _06072_ _06073_ _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10447_ _03194_ _03248_ _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10002__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13166_ _05993_ _06080_ _06082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09943__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10378_ _00517_ _03253_ _03256_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_23_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12117_ _00372_ _00375_ _02236_ _02153_ _04960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_13097_ _05936_ _06007_ _06008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_127_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12048_ _04888_ _04890_ _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_46_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07182__A2 _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09459__A1 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13255__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11266__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08210_ _00989_ _01016_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11018__A1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09190_ _02080_ _02081_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08141_ _01039_ _01042_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09631__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12230__A3 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08072_ _00948_ _00969_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07023_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-10\] _06659_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_151_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08198__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08974_ _00440_ _01782_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07925_ _00823_ _00826_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold49 net19 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XANTENNA__09698__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone7_I net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07856_ _00738_ _00740_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07173__A2 _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07787_ _00709_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06920__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09526_ _02412_ _02413_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09457_ _00357_ _06710_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08408_ _01253_ _01308_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09388_ net61 _06691_ _06696_ net142 _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_81_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08339_ _01215_ _01225_ _01228_ _01229_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_46_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11350_ _04190_ _04191_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10301_ _03003_ _03006_ _03180_ _03172_ _03011_ _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_132_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11980__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11281_ _00372_ _02584_ _02499_ _00375_ _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_131_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13020_ _05861_ _05923_ _05924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10232_ _03049_ _03070_ _03111_ _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11732__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10163_ _00398_ _00394_ _06691_ _06696_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09138__B1 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10094_ _00373_ _06738_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_109_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13922_ _00253_ net36 clknet_leaf_31_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_89_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13853_ _00184_ net36 clknet_leaf_67_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_88_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13237__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12804_ _05687_ _05688_ _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13784_ net126 net36 clknet_leaf_75_clk DDS_Stage.LCU.state\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_10996_ _00381_ _02586_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12735_ _05556_ _05614_ _05615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12666_ _05537_ _05539_ _05541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_13_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11617_ _04287_ _04456_ _04457_ _04458_ _04459_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_115_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12597_ net93 _05462_ _05464_ _05405_ _05428_ _05465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_52_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11548_ _04334_ _04339_ _04390_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11479_ _04218_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13173__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13218_ _06086_ _06101_ _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_133_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13149_ _06056_ _06062_ _06063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07710_ net114 DDS_Stage.xPoints_Generator1.RegF\[-13\] _00667_ _00670_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11487__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08690_ net61 _06649_ _06654_ net60 _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07155__A2 _06732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07641_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-10\] DDS_Stage.xPoints_Generator1.RegFrequency\[-10\]
+ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06902__A2 _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11239__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07572_ _00560_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09311_ _02195_ _02198_ _02201_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_62_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _01982_ _02045_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_32_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_153_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09173_ _01988_ _01989_ _02064_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_145_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08124_ net142 _06179_ _05864_ net61 _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11962__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08055_ _00954_ _00955_ _00956_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_4_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07006_ _06243_ _06623_ _06644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput28 net28 Cos_Out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09907__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11714__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08591__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08957_ _00357_ _06679_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07908_ _00807_ _00808_ _00809_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08888_ _01781_ _01783_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07839_ _00738_ _00739_ _00740_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10150__A1 _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12690__A3 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10850_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[3\] _03674_ _03722_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _02048_ _02145_ _02397_ _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_10781_ _03311_ _03653_ _03585_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08646__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12520_ _03556_ _00354_ _05381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_136_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12451_ _05167_ _05189_ _05308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11402_ _04240_ _04244_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11402__A1 _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12382_ _05211_ _05221_ _05233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11333_ _00387_ _01247_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07082__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07367__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11264_ _00387_ _02153_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13003_ _02938_ _00397_ _05905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10215_ _02929_ _03013_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_11195_ _00397_ _02153_ _03810_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08582__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10146_ _02971_ _02990_ _03026_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13458__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11469__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ _02874_ _02955_ _02958_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07137__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13905_ _00236_ net36 clknet_leaf_23_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_18_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13836_ _00167_ clknet_leaf_71_clk DDS_Stage.xPoints_Generator1.RegP\[-12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10979_ _00361_ _02940_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13767_ _00102_ clknet_leaf_10_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12718_ _05489_ _05499_ _05596_ _05597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13698_ _00033_ clknet_leaf_57_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13870__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12649_ _05516_ _05521_ _05522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_135_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11944__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09860_ _00370_ _06724_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ _01637_ _01651_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_55_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09791_ _02575_ _02666_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08742_ _06637_ _00379_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07128__A2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08673_ _01552_ _01570_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_37_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07624_ DDS_Stage.xPoints_Generator1.CosNew\[-12\] _00597_ _00577_ _00598_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06887__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11880__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07740__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07555_ _05182_ _00548_ _00549_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11632__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11632__B2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07486_ _00492_ _00493_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09225_ net61 net60 _06679_ _06685_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_118_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13861__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09156_ _01967_ _02048_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_5_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08107_ _00997_ _01007_ _01008_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07064__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09087_ _01891_ _01939_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08038_ _00938_ _00939_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_2_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11699__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11699__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ _02704_ _02881_ _02882_ _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09989_ _02779_ _02870_ _02871_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12112__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11951_ _04759_ _04792_ _04793_ _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10902_ _03766_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11882_ _04715_ _04716_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11871__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10833_ _03639_ _03650_ _03638_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13621_ _06571_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10426__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13552_ _06488_ _06497_ _06498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10764_ _03037_ _03579_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_13_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13852__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12503_ _04017_ _04031_ _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13483_ _00384_ _03679_ _06424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10695_ net63 _06742_ net57 _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_109_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__A3 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12179__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12434_ _05283_ _05287_ _05288_ _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07055__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12365_ _05121_ _05122_ _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11316_ _04077_ _04085_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_132_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12296_ net94 _05137_ _05138_ _05140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_50_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11247_ _04087_ _04088_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11178_ _04019_ _04020_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10129_ _02925_ _03010_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_98_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12103__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06869__A1 _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11862__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13819_ _00150_ clknet_leaf_70_clk DDS_Stage.xPoints_Generator1.RegF\[-14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11209__A4 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07340_ _00383_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07294__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07271_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-3\] _00328_ _00329_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11090__A2 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09010_ _01826_ _01902_ _01903_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09035__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11917__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07046__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09912_ _02787_ _02795_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09843_ _02637_ _02638_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10353__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06986_ _05822_ _06627_ _06628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09774_ _02479_ _02483_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08725_ _01548_ _01620_ _01621_ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08849__A2 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ _01397_ _01483_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07607_ _06059_ _00582_ _00583_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08587_ _01406_ _01414_ _01485_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_68_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10408__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11605__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07538_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[0\] _00535_ _00395_ _00536_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10959__A3 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07285__A1 _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07202__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07469_ _06713_ _06211_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ _02026_ _02039_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10480_ _03315_ _03321_ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09139_ net61 net60 _06674_ _06679_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__12030__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12150_ _04990_ _04991_ _04992_ _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11101_ _03939_ _03943_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12081_ _04920_ _04923_ _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_103_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12869__B1 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07645__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11032_ net87 _03340_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10344__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10895__A2 _06765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12983_ _05786_ _05787_ _05883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11934_ _04771_ _04776_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11865_ net66 _01430_ _01249_ net54 _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13604_ _06526_ _06552_ _06553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13597__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10816_ _03401_ _03663_ _03687_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11796_ _04624_ _04637_ _04638_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_144_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07276__A1 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13535_ _06418_ _06428_ _06479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10747_ _03558_ _03620_ _05171_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13466_ _06239_ _06404_ _06406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10678_ _03544_ _03552_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_125_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07028__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12417_ _05262_ _05263_ _05271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13397_ _06330_ _06331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12348_ _04355_ _04409_ _05196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12279_ _04987_ _05005_ _05122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13521__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11678__A4 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ DDS_Stage.LCU.state\[1\] _05226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07200__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08510_ _00357_ _06654_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09490_ _00382_ _06674_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07503__A2 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08441_ _01218_ _01339_ _01340_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13588__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08372_ _01259_ _01272_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_105_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07323_ _00369_ _00370_ _05182_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13816__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07267__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11063__A2 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11602__A4 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07254_ _05182_ _00314_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07019__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07185_ _05452_ _06748_ _06798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07814__I0 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07990__A2 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10326__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_92_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09192__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ _00398_ _06672_ _06674_ _00394_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09731__A3 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12079__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09757_ _02621_ _02642_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06969_ _06059_ _06587_ _06609_ _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08708_ _01533_ _01534_ _01605_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09688_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-11\] _02501_ _02574_ _02575_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_83_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _01535_ _01536_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_25_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13579__A1 _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11650_ _04473_ _04475_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13807__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07258__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10601_ _03405_ _03409_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11581_ _04422_ _04423_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13320_ _06245_ _06246_ _06248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_52_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10532_ _03408_ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_80_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13251_ _06091_ _06100_ _06173_ _06174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_98_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10463_ _05280_ _03340_ _03341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12202_ _05041_ _05044_ _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13182_ _06096_ _06097_ _06098_ _06099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_103_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10394_ _03270_ _03271_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12133_ _04881_ _04885_ _04976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07430__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07375__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07981__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12064_ _04887_ _04905_ _04906_ _04907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _03855_ _03856_ _03857_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12966_ _05759_ _05776_ _05865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_125_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11917_ _00372_ _00375_ _02409_ _02238_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__07497__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13125__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12897_ _05790_ _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11848_ _04656_ _04664_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11779_ _04533_ _04621_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12793__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13518_ _06391_ _06433_ _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_30_clk_I clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13449_ _06333_ _06354_ _06387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08749__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_45_clk_I clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07421__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08990_ _01814_ _01882_ _01883_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_142_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07941_ _06637_ _00355_ _00815_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_103_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07872_ _00773_ _00771_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09713__A3 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[14\] _02499_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_92_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09542_ _02427_ _02428_ _02429_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__11808__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12076__A4 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12481__A1 _05336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09473_ _02360_ _02361_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08424_ _01323_ _01314_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_149_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09229__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ _00916_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12233__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07306_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-13\] _00357_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_73_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08286_ _00951_ _00965_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07237_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-9\] _00301_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12536__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07168_ _05724_ _06629_ _06146_ _06783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07412__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07099_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[1\] _06724_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09809_ net61 _06724_ _06730_ net60 _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12820_ _05608_ _05609_ _05707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_96_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09468__A2 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07479__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11275__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12751_ _05447_ _05537_ _05633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_69_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11702_ net86 _01794_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12682_ _05469_ _05484_ _05557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08691__A3 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11633_ _04474_ _04473_ _04475_ _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_154_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08979__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11564_ _04401_ _04406_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09640__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13303_ _06224_ _06225_ _06228_ _06229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10515_ _03387_ _03391_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11495_ _04336_ _04337_ _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13234_ _06072_ _06073_ _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_122_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10446_ _03269_ _03323_ _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_126_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07403__A1 _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13165_ _05998_ _06080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10377_ _03170_ _03182_ _03255_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10002__A3 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12116_ _04949_ _04952_ _04958_ _04959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13096_ _05938_ _06005_ _06007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_127_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12047_ _00372_ _02238_ _02236_ _00375_ _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07118__B _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_148_Left_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_140_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09459__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11266__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12949_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-9\] _05841_ _05847_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_48_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_72_clk clknet_3_0__leaf_clk clknet_leaf_72_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_105_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12215__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11018__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08140_ _01040_ _01041_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09631__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12230__A4 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08071_ _00971_ _00972_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07022_ _05658_ _06657_ _06658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_141_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08198__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07807__I _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08973_ _01796_ _01798_ _01867_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_07924_ _00824_ _00825_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09698__A2 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07855_ _05833_ _05398_ _00385_ _00382_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_97_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07786_ DDS_Stage.xPoints_Generator1.RegFrequency\[-6\] DDS_Stage.xPoints_Generator1.RegF\[-6\]
+ _00402_ _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09525_ _00370_ _06696_ _02333_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12454__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-23\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_63_clk clknet_3_0__leaf_clk clknet_leaf_63_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09456_ _02281_ _02343_ _02344_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12206__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08407_ _01255_ _01300_ _01307_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_109_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09387_ _02212_ _02216_ _02276_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08338_ _01233_ _01235_ _01239_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10768__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08269_ _06308_ _00370_ _01072_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_62_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10300_ _03171_ _03089_ _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11280_ _00378_ _02409_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10231_ _03030_ _03048_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10162_ _00398_ _06691_ _06696_ _00394_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09138__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09138__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ _02973_ _02974_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07653__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13921_ _00252_ net36 clknet_leaf_31_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_107_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13852_ _00183_ net36 clknet_leaf_69_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__13237__A3 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12803_ _05676_ _05677_ _05686_ _05688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_13783_ _00118_ clknet_leaf_11_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_54_clk clknet_3_1__leaf_clk clknet_leaf_54_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10995_ _00387_ _02499_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12734_ _05591_ _05613_ _05614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_155_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12665_ _05538_ _05448_ _05539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11616_ _04251_ _04252_ _04456_ _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_26_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09613__A2 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12596_ _05391_ _05404_ _05464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11547_ _04329_ _04389_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11478_ _04291_ _04320_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_122_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09377__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13173__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13217_ _03018_ _00397_ _06090_ _06137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_133_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10429_ _00379_ _00376_ _06744_ _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11184__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13148_ _05959_ _06061_ _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10931__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13079_ _03189_ _00390_ _05988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07563__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11487__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07640_ _00611_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07571_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[19\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-12\]
+ _00395_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11239__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09998__B _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_45_clk clknet_3_4__leaf_clk clknet_leaf_45_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09310_ _02199_ _02200_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09241_ _02065_ _02132_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_91_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07863__A1 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09172_ _02063_ _01987_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_153_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08123_ _01023_ _01024_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08054_ net92 net143 _06308_ net153 _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__07738__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07005_ _06059_ _06641_ _06643_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput29 net29 Cos_Out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__11175__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08591__A2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _01758_ _01849_ _01850_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07907_ _00363_ _06627_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08887_ _00440_ _01782_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09540__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08343__A2 _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ _05398_ _00388_ _00385_ _05833_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12690__A4 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07769_ _00700_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_36_clk clknet_3_6__leaf_clk clknet_leaf_36_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09508_ _02396_ _02313_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_10780_ _03388_ _03519_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_137_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09439_ _02258_ _02272_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_109_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12450_ _05297_ _05305_ _05306_ _05307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_81_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11401_ _04241_ _04242_ _04243_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_12381_ _05223_ _05227_ _05232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_133_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11332_ _00390_ _00393_ _01249_ _01247_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__07082__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07209__I1 _06817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11263_ _04072_ _04102_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13002_ _05902_ _05788_ _05903_ _05904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10214_ _03094_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11194_ _03808_ _03809_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10913__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08582__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10145_ _02950_ _02970_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07383__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10076_ net161 _02956_ _02957_ _02779_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11469__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13904_ _00235_ net36 clknet_leaf_20_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_18_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13835_ _00166_ clknet_leaf_71_clk DDS_Stage.xPoints_Generator1.RegP\[-13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_clk clknet_3_7__leaf_clk clknet_leaf_27_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13766_ _00101_ clknet_leaf_10_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10978_ _03817_ _03820_ _03818_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_102_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12717_ _05492_ _05498_ _05596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13697_ _00032_ clknet_leaf_57_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12648_ _05517_ _05519_ _05520_ _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_109_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12579_ _05438_ net145 _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10492__B net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08810_ _01630_ _01683_ _01705_ _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_110_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _01959_ _01966_ _02674_ _02672_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_84_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08741_ _06649_ _00373_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08672_ _01555_ _01569_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07623_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-12\] DDS_Stage.xPoints_Generator1.RegFrequency\[-12\]
+ _00596_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06887__A2 _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11880__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_18_clk clknet_3_7__leaf_clk clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07554_ _00348_ _06733_ _06756_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_49_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07836__A1 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07485_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-10\] _00493_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11632__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone23_I net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09224_ net61 _06679_ _06685_ net60 _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09155_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-17\] _01974_ _02047_ _02048_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_72_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11396__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08106_ net61 net60 _05864_ _05833_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07064__A2 _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09086_ _01887_ _01888_ _01978_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08037_ _00757_ _00759_ _00756_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__11148__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08013__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11699__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09988_ net61 net60 _06738_ _06742_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08939_ _01748_ _01764_ _01833_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_150_Right_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11950_ _04779_ _04791_ _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_4_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10901_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-20\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-20\]
+ _05171_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11881_ _04722_ _04723_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11871__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13620_ net25 _06570_ _05171_ _06571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10832_ _03654_ _03703_ _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_94_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13551_ _06492_ _06496_ _06497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07827__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10763_ _03575_ _03582_ _03635_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12502_ _03979_ _04034_ _05361_ _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13482_ _00387_ _03558_ _06423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10694_ net63 _06742_ net57 _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07842__A4 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12179__A3 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12433_ _05223_ _05227_ _05288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_23_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13620__I0 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11387__A1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07055__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12364_ _05124_ _05212_ _05213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11315_ _04148_ _04156_ _04157_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_112_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12295_ _05135_ _05136_ _05138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_22_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11246_ _04087_ _04088_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09752__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11177_ net135 _00390_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12639__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10128_ _02834_ _02837_ _02924_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10059_ _02916_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11311__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10114__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_121_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06869__A2 _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11862__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13818_ _00149_ clknet_leaf_72_clk DDS_Stage.xPoints_Generator1.RegF\[-15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13064__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07818__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13749_ _00084_ net36 clknet_leaf_48_clk DDS_Stage.xPoints_Generator1.CosNew\[-4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_46_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07270_ _05658_ _00326_ _00327_ _06762_ _05171_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_73_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07294__A2 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09035__A3 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_130_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11917__A3 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07046__A2 _06677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10050__A1 _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09991__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09911_ _02712_ _02794_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09743__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09842_ _02637_ _02638_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10353__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09773_ _02654_ _02658_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06985_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-16\] _06627_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08724_ _01550_ _01599_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08655_ _01479_ _01482_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07606_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-15\] _05280_ _00583_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08586_ _01409_ _01413_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07537_ _00531_ _00532_ _00534_ _05658_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11605__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10959__A4 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08482__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07468_ _00477_ _00478_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09207_ _02026_ _02039_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07399_ _05995_ _00421_ _06254_ _06146_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_20_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09138_ net61 _06674_ _06679_ net60 _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12030__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09069_ _01947_ _01951_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_103_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11100_ _03940_ _03941_ _03942_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__12869__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12080_ _04921_ _04922_ _04805_ _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_112_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12869__B2 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11031_ _00359_ _03189_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10344__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12982_ _05786_ _05787_ _05882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11933_ _04772_ _04775_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_28_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11864_ _04705_ _04706_ _04680_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_156_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13603_ _06529_ _06551_ _06552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10815_ _03082_ _03664_ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13597__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11795_ _04635_ _04636_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13534_ _06473_ _06477_ _06478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_hold86_I FreqPhase[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07276__A2 _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10746_ _03616_ _03619_ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13465_ _06402_ _06403_ _06404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10677_ _03545_ _03547_ _03551_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12416_ _05261_ _05268_ _05270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_23_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13396_ _06320_ _06329_ _06330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_152_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09973__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12347_ _04352_ _05195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12278_ _05108_ _05115_ _05120_ _05121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_121_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13521__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11229_ _04037_ _04038_ _04071_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_52_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07200__A2 _06809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07339__I0 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07571__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_4_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08440_ _01221_ _01222_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13588__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08371_ _01262_ _01266_ _01271_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_59_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07322_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-10\] _00370_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07267__A2 _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06915__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07253_ _05658_ _06623_ _06735_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07184_ _06796_ _06797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07746__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09716__A1 _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07990__A3 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10326__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11523__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09825_ _02708_ _02609_ _02709_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09192__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09731__A4 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13752__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09756_ _02624_ _02627_ _02641_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__12079__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06968_ _05822_ _06598_ _06609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08707_ _01602_ _01604_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_69_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09687_ _02572_ _02573_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06899_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-23\] _05864_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_69_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _01448_ _01449_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08569_ _00388_ _06523_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10600_ _03182_ _03330_ _03474_ _03475_ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_135_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07258__A2 _06623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11580_ _00372_ _01610_ _01524_ _00375_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10531_ _03406_ _03407_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13250_ _06095_ _06172_ _06173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10462_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[24\] _03340_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_114_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12201_ _05042_ _05043_ _05044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10014__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11211__B1 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13181_ _03485_ _00381_ _06098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10393_ _03239_ _03247_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12132_ _04965_ _04973_ _04974_ _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07430__A2 _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12063_ _04903_ _04904_ _04906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11014_ net66 net83 _03189_ _03018_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_95_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13743__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06941__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07391__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12965_ _05794_ _05817_ _05862_ _05863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_125_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11916_ _04747_ _04752_ _04758_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08694__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12896_ _05784_ _05788_ _05790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11847_ _04679_ _04688_ _04689_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_51_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11778_ _04531_ _04532_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13517_ _06393_ _06432_ _06460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10729_ _03602_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13448_ _06335_ _06353_ _06386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08749__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09946__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13379_ _06262_ _06280_ _06312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07957__B1 _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07421__A2 _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07940_ _00788_ _00818_ _00841_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07871_ _00772_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09713__A4 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07185__A1 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13734__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09610_ _02496_ _02497_ _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06932__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09541_ net142 _06710_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11808__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09472_ _06654_ _00394_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10492__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08423_ _00980_ _00930_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08354_ _00907_ _00925_ _01254_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12233__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10244__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07305_ _00356_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08285_ _01053_ _01089_ _01186_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_rebuffer33_I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06999__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07236_ _06624_ _00299_ _05658_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07167_ _05387_ _06777_ _06782_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07412__A2 _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07098_ _06146_ _06722_ _06723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_93_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13725__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09808_ _02605_ net149 _02692_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06923__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09739_ _02533_ _02536_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12750_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-11\] _05631_ _05632_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11701_ _04541_ _04542_ _04543_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11680__B1 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12681_ _05502_ _05524_ _05555_ _05556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08691__A4 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11632_ _00361_ _01792_ _01693_ _00365_ _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10235__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11563_ _04402_ _04405_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07100__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13302_ _06174_ _06226_ _06227_ _06228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10514_ _03388_ _03389_ _03390_ _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_24_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11494_ _00390_ _01430_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13233_ _06150_ _06153_ _06154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_134_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09928__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10445_ _03272_ _03322_ _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13164_ _06055_ _06078_ _06079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_hold49_I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07403__A2 _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10376_ _03166_ _03254_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10002__A4 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12115_ _04953_ _04957_ _04958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13095_ _06004_ _06005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09156__A2 _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12046_ _00378_ _02153_ _04889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07167__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06914__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08667__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12948_ _05732_ _05846_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13660__A1 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11266__A3 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12879_ _03556_ _00369_ _05771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13412__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12215__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09631__A3 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11974__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08070_ _00770_ _00820_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07021_ _06615_ _06656_ _06657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13955__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08972_ _01863_ _01866_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07923_ net155 _00376_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07158__A1 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12151__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07854_ _00750_ _00755_ _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10162__B1 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06905__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07785_ _00708_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clone53_I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09524_ _02411_ _02332_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08658__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09455_ net91 net142 _06696_ _06701_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_149_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08406_ _01301_ _01306_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_35_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13403__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12206__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09386_ _02207_ _02211_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08337_ _01236_ _01238_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11414__B1 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10768__A2 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08268_ _00984_ _01095_ _01169_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_117_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07219_ _05669_ _06688_ _06826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ _01099_ _01100_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_132_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10230_ _03108_ _03109_ _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07397__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13946__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10161_ _02704_ _03040_ _03041_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09138__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10092_ _02792_ _02887_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07149__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13920_ _00251_ net36 clknet_leaf_32_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_22_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08897__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13851_ _00182_ net36 clknet_leaf_72_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_69_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12802_ _05676_ _05677_ _05686_ _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_122_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13782_ _00117_ clknet_leaf_4_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08649__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10994_ _03802_ _03836_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12733_ _05595_ _05597_ _05612_ _05613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA_clkbuf_leaf_44_clk_I clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12664_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-13\] _05446_ _05538_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11615_ _04420_ _04435_ _04437_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_143_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09074__A1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12595_ _05391_ _05404_ _05462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_80_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_59_clk_I clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11546_ _04333_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_123_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11477_ _04307_ _04319_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13216_ _06088_ _06089_ _06136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10428_ _03301_ _03305_ _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09377__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13937__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11184__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13147_ _06057_ _06060_ _06061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10359_ _03214_ _03237_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13078_ _03018_ _00393_ _05987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12029_ _04800_ _04861_ _04871_ _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__10695__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07560__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07570_ _00559_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09240_ _02068_ _02131_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_119_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07863__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09171_ _01985_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08122_ _01021_ _01022_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08053_ net92 _06308_ _06416_ _00363_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07004_ _05822_ _06642_ _06643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13928__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11175__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07754__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08955_ net61 net142 _06664_ _06672_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_110_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12124__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07906_ _00367_ _06618_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08886_ _01775_ _01780_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10686__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09540__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07837_ _05864_ _00382_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_16_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07551__A1 _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_1__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07768_ DDS_Stage.xPoints_Generator1.RegFrequency\[-15\] DDS_Stage.xPoints_Generator1.RegF\[-15\]
+ _00402_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09507_ _00463_ _02156_ _02227_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_94_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _00660_ _00661_ _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09438_ _02251_ _02303_ _02326_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09369_ _00373_ _06685_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11400_ _00359_ _02153_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_25_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07606__A2 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12380_ _05211_ _05221_ _05231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11331_ _04106_ _04173_ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__10610__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11262_ _04036_ _04104_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13919__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13001_ _05781_ _05791_ _05903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10213_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-5\] _03091_ _03093_ _03094_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_123_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11193_ _03850_ _03971_ _04035_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__10913__A2 _06811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08582__A3 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10144_ _03023_ _03024_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10075_ _02873_ _02874_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_34_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11469__A3 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13903_ _00234_ net36 clknet_leaf_20_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07542__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13834_ _00165_ clknet_leaf_70_clk DDS_Stage.xPoints_Generator1.RegP\[-14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10429__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11626__B1 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13765_ _00100_ clknet_leaf_9_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10977_ _03818_ _03819_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09295__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12716_ _05513_ _05522_ _05593_ _05595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13696_ _00031_ clknet_leaf_54_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12647_ _02940_ _00381_ _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_135_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12578_ _05250_ _05270_ _05439_ _05444_ _05445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_29_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11529_ _04316_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08740_ _01635_ _01636_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08671_ _01560_ _01568_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11865__B1 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07533__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07622_ _00594_ _00595_ _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07553_ _06092_ _06622_ _00547_ _05658_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_48_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07836__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07484_ _05182_ _00490_ _00491_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_124_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09223_ _02112_ _02113_ _02114_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09038__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09154_ _02046_ _01976_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08105_ net60 _05864_ _05833_ net61 _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11396__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09085_ _01977_ _01886_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08036_ _00933_ _00937_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11148__A2 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08013__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10903__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09987_ net61 _06738_ _06742_ net60 _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08938_ _01750_ _01763_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10659__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08869_ _01748_ _01764_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10900_ _05822_ _06777_ _03765_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_4_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11880_ _00361_ _01247_ _04713_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10831_ _03592_ _03702_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13550_ _06493_ _06494_ _06495_ _06496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_39_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10762_ _03577_ _03580_ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12501_ _03981_ _04033_ _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13481_ _06421_ _06422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10693_ _03505_ _03511_ _03566_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12432_ _04742_ _05284_ _05285_ _05286_ _05287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07659__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12179__A4 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13620__I1 _06570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11387__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12363_ _05127_ _05212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_121_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11314_ _04152_ net81 _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12294_ _05135_ _05136_ _05137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_130_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11245_ _03863_ _03864_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09201__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10898__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09752__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11176_ _00393_ _02499_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10127_ _03008_ _02926_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12639__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[20\] _02940_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_54_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11311__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13817_ _00148_ net36 clknet_leaf_46_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__13064__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07818__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13748_ _00083_ net36 clknet_leaf_48_clk DDS_Stage.xPoints_Generator1.CosNew\[-5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_45_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13679_ _00014_ clknet_leaf_0_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_42_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07569__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09035__A4 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11917__A4 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09991__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09910_ _02790_ _02793_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09841_ _02722_ _02725_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_70_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09743__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09772_ _02655_ _02657_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06984_ _06146_ _06625_ _06626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08723_ _01550_ _01599_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11838__B1 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07506__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08654_ _01463_ _01471_ _01551_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_1_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07605_ DDS_Stage.xPoints_Generator1.CosNew\[-15\] _00578_ _00579_ _00581_ _00582_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_139_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08585_ _01397_ _01483_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09259__A1 _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07536_ _06232_ _05919_ _00533_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07467_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-13\] _00478_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08482__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09206_ _02079_ _02097_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_17_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07398_ _05409_ _05897_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09137_ _02027_ _02028_ _02029_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_103_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09068_ _01775_ _01949_ _01960_ _01950_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07442__B1 _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08019_ _00919_ _00920_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10329__B1 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12869__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11030_ _03859_ _03871_ _03872_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_9_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12981_ _05869_ _05880_ _05881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11932_ _04773_ _04774_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_59_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11863_ net54 _01430_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_28_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10814_ _03629_ _03684_ _03685_ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_13602_ _06532_ _06533_ _06550_ _06551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_67_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11057__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13597__A3 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11794_ _04635_ _04636_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_156_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13533_ _06239_ _06476_ _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_137_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10745_ _03618_ _03554_ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07389__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13464_ _06323_ _06396_ _06401_ _06403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10676_ _03549_ _03550_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_153_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12557__A1 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12415_ _05264_ _05267_ _05268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_3_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13395_ _06239_ _06328_ _06329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12346_ _04348_ _04351_ _05194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_2_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12277_ _05106_ _05107_ _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11228_ _04051_ _04069_ _04070_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07736__A1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11159_ _03934_ _03935_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07339__I1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11048__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08370_ _01267_ _01270_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07321_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-10\] _00369_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_46_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09661__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07252_ _06232_ _06351_ _06681_ _05550_ _05658_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_73_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_143_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12548__A1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07183_ _05507_ _06795_ _05647_ _06796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09716__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07990__A4 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11523__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12720__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09824_ net63 _06674_ _02608_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07762__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06967_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-18\] _06598_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09755_ _02632_ _02640_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08706_ _01440_ _01505_ _01603_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11287__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09686_ _02502_ _02503_ _02571_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06898_ _05811_ _05844_ _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08637_ _01445_ _01446_ _01444_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_25_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08568_ _00382_ _06618_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12787__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07519_ _05658_ _06623_ _00465_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08499_ _01371_ _01395_ _01398_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_37_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10530_ _03269_ _03323_ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10461_ _03336_ _03338_ _03339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12200_ _00372_ _02153_ _02051_ _00375_ _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11211__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10014__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13180_ net147 _00384_ _06097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10392_ _03196_ _03238_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11211__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12131_ _04971_ _04972_ _04974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12062_ _04903_ _04904_ _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07569__I1 DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_11013_ net66 _03189_ _03018_ net83 _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_8_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06941__A2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12964_ _05757_ _05793_ _05862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_125_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11915_ _04753_ _04757_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12895_ _05785_ _05786_ _05787_ _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08694__A2 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11846_ _04683_ _04687_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11777_ _04615_ _04619_ _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10728_ _03596_ _03601_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13516_ _06388_ _06390_ _06459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_83_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10659_ _03082_ _03533_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13447_ _06382_ _06357_ _06384_ _06385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09946__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13378_ _06262_ _06280_ _06311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07957__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07957__B2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12329_ _05170_ _05174_ _05175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07870_ net58 _06633_ _06627_ _00355_ _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08382__A1 _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06932__A2 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09540_ net92 _06708_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11269__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09471_ _06649_ _00398_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08422_ _01312_ _01321_ _01310_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_TAPCELL_ROW_65_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10492__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout36_I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08353_ _00880_ _00906_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09634__A1 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07304_ net54 _00355_ _05182_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08284_ _01087_ _01088_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07235_ _05409_ _06211_ _06756_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07166_ _06146_ _06778_ _06781_ _05182_ _06782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07948__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07097_ _06720_ _06721_ _06722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_140_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09807_ net150 _02604_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13507__B DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07999_ _06654_ _00352_ _00391_ _05864_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06923__A2 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09738_ _02550_ _02558_ _02623_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08125__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09873__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09669_ _00385_ _06679_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11700_ net66 net54 _01792_ _01693_ _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07884__B1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11680__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12680_ _05466_ _05462_ _05501_ _05555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11680__B2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11631_ _00369_ _01610_ _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_145_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10235__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11562_ _04403_ _04404_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_53_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07100__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10513_ _00385_ _06742_ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13301_ _06177_ _06193_ _06227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_108_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11493_ _00393_ _01249_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13232_ _05959_ _06152_ _06153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07667__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10444_ _03315_ _03321_ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09928__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_clk_I clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13163_ _06063_ _06077_ _06078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10375_ _03169_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12114_ _04954_ _04955_ _04956_ _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_130_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13094_ _05946_ _06003_ _06004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12045_ _00372_ _00375_ _02238_ _02236_ _04888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_127_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07167__A2 _06777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08364__A1 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12947_ _05387_ _05843_ _05845_ _05846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08667__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13660__A2 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11266__A4 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12878_ _05763_ _05769_ _05770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_47_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11829_ _04670_ _04671_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_145_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13412__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11423__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07150__B _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10226__A2 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_155_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09631__A4 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11974__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07577__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07020_ _05409_ _05940_ _06656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08971_ _01704_ _01864_ _01865_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_07922_ net152 _00379_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12151__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ _00753_ _00754_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10162__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10162__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07784_ DDS_Stage.xPoints_Generator1.RegFrequency\[-7\] DDS_Stage.xPoints_Generator1.RegF\[-7\]
+ _00402_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09523_ _02330_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08658__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09454_ net91 _06696_ _06701_ net142 _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08405_ _01303_ _01305_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_149_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13891__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09385_ _02202_ _02218_ _02274_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_35_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13403__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12206__A3 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08336_ _00984_ net71 _01237_ _01169_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__11414__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11414__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10768__A3 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08267_ _01069_ _01094_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_62_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07218_ _05409_ _05550_ _06092_ _06622_ _05658_ _06825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_TAPCELL_ROW_95_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08198_ _00355_ _06179_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_89_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _06146_ _06716_ _06766_ _06767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_30_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10160_ net63 _06696_ _02608_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13946__CLK clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10091_ _02883_ _02886_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08346__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10153__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08897__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13850_ _00181_ net36 clknet_leaf_71_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_98_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12801_ _05681_ _05685_ _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13781_ _00116_ clknet_leaf_4_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08649__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10993_ _03802_ _03801_ _03803_ _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09846__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12732_ _05602_ _05611_ _05612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13882__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12663_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-12\] _05536_ _05537_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11614_ _04251_ _04252_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_13_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11405__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12602__B1 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09074__A2 _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12594_ _05458_ _05460_ _05461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_80_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07085__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_137_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11545_ _04371_ _04385_ _04387_ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_107_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13158__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold61_I FreqPhase[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11476_ _04310_ _04318_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ _03302_ _03303_ _03304_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_13215_ _06050_ _06105_ _06133_ _06134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_150_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13146_ _05957_ _06058_ _06060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_10358_ _03218_ _03221_ _03236_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_13077_ _02940_ _00397_ _05986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10289_ _03022_ _03167_ _03168_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_100_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12028_ _04863_ _04864_ _04870_ _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_73_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10695__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07560__A2 _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09837__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11644__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13873__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09170_ _02060_ _02061_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_16_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08121_ _01021_ _01022_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07076__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08052_ net73 _06523_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07003_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-13\] _06642_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_142_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11580__B1 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08954_ net61 _06664_ _06672_ net142 _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12124__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07905_ _00357_ _06633_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08885_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-20\] _01775_ _01780_ _01781_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__07000__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07836_ _05833_ _05398_ _00388_ _00385_ _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__07770__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07767_ _00699_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09506_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-13\] _02394_ _02395_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_79_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07698_ DDS_Stage.xPoints_Generator1.RegFrequency\[-2\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-2\]
+ _00656_ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13864__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09437_ _02253_ _02302_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13388__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09368_ _02195_ _02256_ _02257_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08319_ _01206_ _01210_ _01220_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_118_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09299_ _02185_ _02189_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11330_ _04141_ _04145_ _04172_ _04171_ _04170_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__10610__A2 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11261_ _04072_ _04102_ _04103_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_132_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13000_ _05784_ _05902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10212_ _03007_ _03012_ _03092_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_132_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11192_ _03979_ _04034_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10143_ _02992_ _03000_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08582__A4 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13312__A1 _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10074_ _02873_ _02874_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11469__A4 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13902_ _00233_ net36 clknet_leaf_21_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07680__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07542__A2 _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13833_ _00164_ clknet_leaf_73_clk DDS_Stage.xPoints_Generator1.RegP\[-15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10429__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11626__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11626__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13764_ _00099_ clknet_leaf_1_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10976_ _00372_ _02762_ _02586_ _00375_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09295__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13855__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12715_ _05516_ _05592_ _05593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13695_ _00030_ clknet_leaf_6_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12646_ _02938_ _00384_ _05519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07058__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12051__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12577_ _05443_ _05444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11528_ _04357_ _04370_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_29_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11459_ _00369_ _02051_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07230__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13129_ _05948_ _06002_ _06042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10117__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08670_ _01563_ _01567_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11865__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11865__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07533__A2 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07621_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\] DDS_Stage.xPoints_Generator1.RegFrequency\[-13\]
+ _00590_ _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07552_ _05550_ _06789_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07297__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07483_ _05658_ _05529_ _06651_ _06712_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_124_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07836__A3 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09222_ net58 _06708_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09038__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07049__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09153_ _01979_ _01982_ _02045_ _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_146_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08104_ _01004_ _01005_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_12_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08797__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11396__A3 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09084_ _01884_ _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08035_ _00934_ _00935_ _00936_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_141_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_43_clk_I clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09986_ _02783_ _02785_ _02868_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08937_ _01814_ _01817_ _01831_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_08868_ _01750_ _01763_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_clkbuf_leaf_58_clk_I clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07819_ _06059_ _00567_ _00725_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08799_ _01530_ _01605_ _01531_ _01687_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_10830_ _03700_ _03701_ _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07288__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10761_ _03584_ _03594_ _03633_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12500_ _05326_ _05355_ _05357_ _05358_ _05359_ _05360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_10692_ _03507_ _03510_ _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13480_ _06347_ _06419_ _06420_ _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12431_ _05245_ _05246_ _05286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_124_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08344__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12362_ _04985_ _05210_ _05211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_50_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11313_ _04152_ _04155_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07460__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12293_ _05026_ _05031_ _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_132_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13533__A1 _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11244_ _04077_ _04085_ _04086_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09201__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07212__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11175_ _00397_ _02409_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10898__A2 _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10126_ _02838_ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10057_ _02935_ _02937_ _02939_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13816_ _00147_ net36 clknet_leaf_45_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_86_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07279__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13747_ _00082_ net36 clknet_leaf_49_clk DDS_Stage.xPoints_Generator1.CosNew\[-6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10959_ _00381_ _00384_ _02584_ _02499_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_128_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13678_ _00013_ clknet_leaf_77_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12629_ _05489_ _05499_ _05500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08779__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11783__B1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07451__A1 _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07451__B2 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07203__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09840_ _02723_ _02724_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08951__A1 _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09771_ _02506_ _02655_ _02656_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06983_ _06620_ _06622_ _06623_ _06624_ _06625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08722_ _01617_ _01618_ _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11838__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11838__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08653_ _01466_ _01470_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07604_ _00578_ _00580_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08584_ _01479_ _01482_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_85_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07535_ _06645_ _06748_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ _00473_ _00474_ _00476_ _05658_ _05182_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_147_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10694__B net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09205_ _02082_ _02096_ _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ _05658_ _06779_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09136_ _06637_ net95 _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10577__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07442__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09067_ _01947_ _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07993__A2 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08018_ _06598_ _00376_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10329__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10329__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07508__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09969_ _02850_ _02852_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12980_ _05873_ _05879_ _05880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11931_ _00372_ _02499_ _02409_ _00375_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11862_ net66 _01524_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13601_ _06539_ _06549_ _06550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10813_ _03632_ _03666_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11057__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11793_ _04549_ _04551_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13532_ _06474_ _06475_ _06476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10744_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[1\] _03617_ _03618_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13463_ _06323_ _06396_ _06401_ _06402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10675_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-1\] _03482_ _03548_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[0\]
+ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_36_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07808__I0 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12414_ _04800_ _05265_ _05266_ _05267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12557__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13394_ _06321_ _06327_ _06328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_23_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12345_ _05176_ _05185_ _05186_ _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_121_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12276_ _05069_ _05117_ _05118_ _05119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_120_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11227_ _04067_ _04068_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_120_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_147_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08933__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11158_ _03934_ _03935_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10109_ _02971_ _02990_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11089_ _03902_ _03910_ _03931_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11048__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07320_ _00368_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09661__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07251_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-6\] _00312_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_45_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12548__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ _05409_ _05529_ _06795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10559__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_52_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08924__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09823_ net63 _06674_ _02608_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12720__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09754_ _02635_ _02639_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06966_ _05658_ _06576_ _06587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08705_ _01442_ _01504_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11287__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_61_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09685_ _02502_ _02503_ _02571_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06897_ _05822_ _05833_ _05844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10495__B1 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08636_ _01328_ _01348_ _01432_ _01508_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_139_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12236__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08567_ _01382_ _01464_ _01465_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12787__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07518_ _05713_ _06614_ _00518_ _05658_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08498_ _01396_ _01397_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_76_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_147_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07449_ _05387_ _00459_ _00460_ _00462_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_119_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10460_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-3\] _03337_ _03263_ _03338_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_70_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_98_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07415__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09119_ _01997_ _02011_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11211__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07415__B2 _06732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10391_ _03242_ _03245_ _03268_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12130_ _04971_ _04972_ _04973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_102_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12061_ _04753_ _04757_ _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11012_ _00359_ _02940_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12963_ _05857_ _05860_ _05861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08679__B1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11914_ _04754_ _04755_ _04756_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_59_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12894_ _03485_ _00372_ _05787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11845_ _04683_ _04687_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11776_ _04617_ _04618_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_126_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13515_ _06455_ _06456_ _06457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10727_ _03082_ _03600_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_153_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13446_ _06318_ _06356_ _06384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10658_ _03401_ _03532_ _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_141_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07406__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13377_ _03266_ _00397_ _06267_ _06310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10589_ _03082_ _03464_ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_106_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07957__A2 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12328_ _05173_ _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12259_ _05034_ _05061_ _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_103_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08382__A2 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11269__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_75_clk clknet_3_0__leaf_clk clknet_leaf_75_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_116_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09470_ _02286_ _02357_ _02358_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08421_ _00767_ _00929_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07893__A1 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_127_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07611__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08352_ _00876_ _00927_ _01252_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09634__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11977__B1 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07303_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-14\] _00355_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
XFILLER_0_156_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08283_ _01184_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07234_ _06211_ _06687_ _06146_ _06006_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09398__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07165_ _05431_ _06779_ _06780_ _06781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07948__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07096_ _05420_ _05886_ _06232_ _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__10952__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_136_Left_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_93_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10704__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11901__B1 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09806_ net151 _02611_ _02688_ _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_07998_ _06654_ _00352_ _00391_ _05864_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__12457__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-21\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09737_ _02553_ _02622_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06949_ _06146_ _06394_ _06405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08125__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_66_clk clknet_3_1__leaf_clk clknet_leaf_66_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09322__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09668_ _00388_ _06674_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12209__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08619_ _01515_ _01516_ _01517_ _01511_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07884__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07884__B2 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11680__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09599_ _02310_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_11630_ _00361_ _00365_ _01792_ _01693_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_49_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11561_ _00390_ _01524_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13300_ _06177_ _06193_ _06226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10512_ _00388_ _06738_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11492_ _00397_ _01247_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09389__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13231_ _06060_ _06151_ _06152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10443_ _03082_ _03320_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11196__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13162_ _06066_ _06076_ _06077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10374_ _03249_ _03252_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12113_ _00393_ _01693_ _04956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13093_ _05948_ _06002_ _06003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_20_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12044_ _04877_ _04880_ _04886_ _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12696__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08364__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12448__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-24\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_clk clknet_3_3__leaf_clk clknet_leaf_57_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12946_ _05740_ _05842_ _05845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11120__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07875__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12877_ _05766_ _05768_ _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_75_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11828_ _04635_ _04636_ _04624_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_28_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11423__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11759_ _04594_ _04595_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_154_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13429_ _06210_ _06294_ _06366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08052__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08970_ _01706_ _01769_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07921_ _06598_ _00373_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12687__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07852_ _00751_ _00752_ _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10162__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12439__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 net134 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07783_ _00707_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_48_clk clknet_3_4__leaf_clk clknet_leaf_48_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09522_ _02406_ _02408_ _02410_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09453_ _02285_ _02289_ _02341_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08404_ _00918_ _00921_ _01304_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_clone39_I net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09384_ _02204_ _02217_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_35_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12206__A4 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08335_ _01195_ _01173_ _01192_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__12611__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11414__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07768__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08266_ _01096_ _01167_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08418__I0 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07217_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-12\] _06824_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_95_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08197_ net58 _06308_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_144_Left_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_131_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07148_ _06447_ _06688_ _06766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07079_ _05930_ _06705_ _06706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10090_ _02900_ _02909_ _02907_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08346__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10153__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_39_clk clknet_3_5__leaf_clk clknet_leaf_39_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12800_ _05682_ _05683_ _05684_ _05685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_153_Left_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13780_ _00115_ clknet_leaf_5_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10992_ _03821_ _03833_ _03834_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_122_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09846__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12731_ _05606_ _05610_ _05611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_139_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12662_ _05530_ _05532_ _05535_ _05536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_93_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11613_ _04441_ _04454_ _04455_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__12602__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11405__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12602__B2 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12593_ _05413_ _05414_ _05459_ _05460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11544_ _04307_ _04319_ _04386_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_80_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13158__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11475_ _04313_ _04317_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_21_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13214_ _06052_ _06104_ _06133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10426_ _00385_ _06738_ _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08034__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10916__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13145_ _00365_ _03727_ _06058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10357_ _03227_ _03235_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13076_ _05982_ _05892_ _05983_ _05985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12669__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10288_ _03025_ _03084_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_12027_ _04866_ _04869_ _04870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07426__B _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10695__A3 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09837__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07848__A1 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12929_ _05643_ _05719_ _05826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11644__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08120_ _00355_ net155 _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07076__A2 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10080__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08051_ _00952_ _00951_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_43_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07002_ _06639_ _06640_ _06641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_77_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10907__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11580__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11580__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08953_ _01845_ _01846_ _01847_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_110_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09525__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07904_ _00793_ _00804_ _00805_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08884_ _01776_ _01778_ _01779_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11332__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07835_ _00730_ _00735_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07000__A2 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13085__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07766_ net7 DDS_Stage.xPoints_Generator1.RegP\[-1\] _00684_ _00699_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_2_clk_I clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09505_ _02319_ _02393_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07697_ DDS_Stage.xPoints_Generator1.RegFrequency\[-2\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-2\]
+ _00660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09436_ _02323_ _02324_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13388__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09367_ _02198_ _02201_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10917__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11399__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08318_ _01208_ _01209_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09298_ _02186_ _02187_ _02188_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_117_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10071__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08249_ _01149_ _01150_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_119_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08016__A1 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11260_ _04100_ _04101_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10211_ _03003_ _03006_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_132_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11191_ _03981_ _04033_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11571__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10142_ _02947_ _02991_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10073_ net61 _06744_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07246__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13901_ _00232_ net36 clknet_leaf_22_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_13832_ _00163_ clknet_leaf_43_clk DDS_Stage.xPoints_Generator1.RegF\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13763_ _00098_ clknet_leaf_12_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12823__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11626__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10975_ _00372_ _00375_ _02762_ _02586_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_12714_ _05521_ _05592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_44_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13694_ _00029_ clknet_leaf_6_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12645_ _02854_ _00387_ _05517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07058__A2 _06125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12051__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12576_ _04036_ _04104_ _05275_ _05439_ _05441_ _05443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_81_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_152_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11527_ _04369_ _04365_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11458_ _04296_ _04300_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_21_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10409_ _00398_ _00394_ _06708_ _06710_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_68_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11389_ net70 _02051_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13128_ _05943_ _05944_ _05942_ _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13791__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13059_ _05871_ _05872_ _05966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_139_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10117__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11865__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\] DDS_Stage.xPoints_Generator1.RegFrequency\[-13\]
+ _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07533__A3 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07551_ _00545_ _00546_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12814__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07482_ _00450_ _00489_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07836__A4 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09221_ _06642_ net98 _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09152_ _02044_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_133_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08103_ net58 _00355_ net152 net155 _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_114_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09994__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08797__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11396__A4 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09083_ _01878_ _01942_ _01975_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_142_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08034_ _05864_ _00379_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09985_ _02778_ _02782_ _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08936_ _01822_ _01830_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_122_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06980__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08867_ _01754_ _01762_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07818_ _05280_ _00385_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08798_ _06059_ _01692_ _01694_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07749_ _00690_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10220__B _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10760_ _03567_ _03583_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09419_ _02161_ _02307_ _02308_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10691_ _03513_ _03527_ _03564_ _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12430_ _05164_ _05190_ _05242_ _05243_ _05285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__13230__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12361_ _05011_ _05012_ _05210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11312_ _04153_ _04154_ _04078_ _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_12292_ _04375_ _04384_ _05134_ _05135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11243_ _04081_ _04084_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11174_ _03919_ _03929_ _04016_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10125_ _03003_ _03006_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__06971__A1 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10056_ _05280_ _02938_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13049__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13815_ _00146_ net36 clknet_leaf_46_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13746_ _00081_ net36 clknet_leaf_51_clk DDS_Stage.xPoints_Generator1.CosNew\[-7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08476__A1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10958_ _00387_ _02409_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10283__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13677_ _00012_ clknet_leaf_77_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10889_ _03759_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12628_ _05492_ _05498_ _05499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_42_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08779__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09976__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12559_ _05421_ _05422_ _05423_ _05424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__11783__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11783__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08400__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07203__A2 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08951__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09770_ _02509_ _02570_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06982_ _06232_ _06620_ _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__13288__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06962__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08721_ _01546_ _01547_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11838__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09900__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ _01474_ _01502_ _01549_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_1_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07603_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-15\] DDS_Stage.xPoints_Generator1.RegFrequency\[-15\]
+ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08583_ _01480_ _01481_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07534_ _06232_ _05897_ _05658_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13460__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07465_ _05442_ _00475_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clone21_I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ _02087_ _02095_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_rebuffer49_I _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13212__A1 _05740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07396_ _05409_ _06714_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_45_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09135_ net58 _06701_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10577__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09066_ _01788_ _01784_ _01958_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_60_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08017_ net156 _00379_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10329__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09968_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-9\] _02851_ _02760_ _02852_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06953__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08919_ _01726_ _01734_ _01813_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09899_ _02778_ _02782_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10888__I0 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11930_ _00372_ _00375_ _02499_ _02409_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__07902__B1 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11861_ _04645_ _04674_ _04697_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_68_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13600_ _06543_ _06548_ _06549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10812_ _03632_ _03666_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_28_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13451__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11792_ _04632_ _04633_ _04634_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_94_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13531_ _06323_ _06398_ _06401_ _06475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_10743_ _03613_ _03543_ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07130__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13462_ _06244_ _06400_ _06401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13203__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10674_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[0\] _03548_ _03549_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_153_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12413_ _04861_ _04871_ _05266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13393_ _06244_ _06326_ _06327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_129_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12344_ _05164_ _05190_ _05191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_51_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__A1 _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12275_ _05104_ _05116_ _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11226_ _04067_ _04068_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13746__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07197__B2 _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08933__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11157_ _03924_ _03927_ _03925_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_52_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06944__A1 _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10108_ _02972_ _02975_ _02989_ _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_65_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11088_ _03905_ _03909_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10039_ _02913_ _02921_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08449__A1 _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11048__A3 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_42_clk_I clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13729_ _00064_ net36 clknet_leaf_16_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_14_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07121__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07250_ _00311_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09949__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07181_ _06793_ _06794_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_57_clk_I clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13737__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09822_ _02693_ _02706_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_6_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08924__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06935__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09753_ _02636_ _02637_ _02638_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06965_ _05409_ _06081_ _06555_ _06566_ _05431_ _06576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_08704_ _01537_ _01601_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08688__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09684_ _02506_ _02509_ _02570_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06896_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-24\] _05833_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10495__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08635_ _01532_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10495__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08566_ _01383_ _01384_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_25_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12236__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13433__A1 _06131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ _05875_ _06666_ _06613_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _06179_ _00398_ _05864_ _00394_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_71_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07112__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07448_ _05182_ _00461_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08860__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07379_ DDS_Stage.xPoints_Generator1.CosNew\[-8\] DDS_Stage.xPoints_Generator1.RegP\[-8\]
+ _00402_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10925__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09118_ _02002_ _02010_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_98_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10390_ _03082_ _03246_ _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09049_ _01878_ _01942_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12060_ _04893_ _04901_ _04902_ _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07179__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13728__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11011_ _03821_ _03833_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06926__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08679__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12962_ _05858_ _05859_ _05860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08679__B2 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10486__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11913_ _00393_ _01794_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12893_ net147 _00375_ _05786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13900__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11844_ _04684_ _04685_ _04686_ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_32_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10238__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11775_ _00369_ _01249_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07103__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold84_I FreqPhase[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10726_ _03401_ _03599_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13514_ _06314_ _06435_ _06456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13445_ _06316_ _06382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10657_ _03446_ _03530_ _03531_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_70_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13376_ _06264_ _06266_ _06309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10588_ _03401_ _03463_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_140_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12327_ _04403_ _04404_ _05172_ _05173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07429__B _06646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09159__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12258_ _05087_ _05100_ _05101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_142_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11209_ _00372_ _00375_ _02586_ _02584_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_103_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12189_ _05025_ _05032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07590__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07164__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13663__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11269__A3 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10477__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07193__I1 _06804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08420_ _00418_ _01317_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_116_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_82_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07893__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08351_ _00878_ _00926_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_46_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11977__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07302_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-14\] _00354_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_156_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11977__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08282_ _01182_ _01183_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07233_ _05387_ _00296_ _00297_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09398__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07164_ _06232_ _06644_ _05658_ _06780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_30_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10401__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07948__A3 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07095_ _05420_ _06092_ _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10952__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_93_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06908__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10704__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11901__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11901__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _02595_ _02688_ _02689_ _02621_ _02642_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_07997_ _06649_ _00355_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06948_ _06362_ _06383_ _06394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09736_ _02557_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08125__A3 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09322__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09667_ _00382_ _06685_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06879_ DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[4\] _05647_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_96_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08618_ _01346_ _01230_ _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_139_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07884__A2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12209__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09598_ _02484_ _02485_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08549_ _01447_ _01444_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11968__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11560_ _00393_ _01430_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10235__A4 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10511_ _00382_ _06744_ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10640__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11491_ _04329_ _04333_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13230_ _00369_ _03727_ _06151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10442_ _03318_ _03319_ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09389__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13949__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11196__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08597__B1 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13161_ _06075_ _06076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_131_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10373_ _03250_ _03251_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12112_ _00390_ _01792_ _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13092_ _05978_ _06001_ _06002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12043_ _04881_ _04885_ _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12696__A2 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12945_ _05740_ _05842_ _05843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11120__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12876_ net70 _03725_ _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07875__A2 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11827_ _04654_ _04668_ _04669_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11758_ _04416_ _04589_ _04590_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10709_ _03575_ _03582_ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10631__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11689_ _00375_ _01247_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13428_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-3\] _06364_ _06365_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_51_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12384__A1 _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08588__B1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13359_ _06200_ _06203_ _06291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08052__A2 _06523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07920_ _00770_ _00820_ _00821_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12687__A2 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10698__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ _00751_ _00752_ _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_78_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08760__B1 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 net122 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07782_ DDS_Stage.xPoints_Generator1.RegFrequency\[-8\] DDS_Stage.xPoints_Generator1.RegF\[-8\]
+ _00402_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13636__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12439__A2 _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09521_ _05280_ _02409_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09452_ _02280_ _02284_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08403_ _00919_ _00920_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09383_ _02255_ _02258_ _02272_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10539__I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[25\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08334_ _01195_ _01193_ _01235_ _01196_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_47_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12611__A2 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08265_ _01119_ _01120_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07216_ _06823_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08196_ _05398_ _00373_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-23\] _06765_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07784__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07078_ _06703_ _06704_ _06705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09719_ _02600_ _02604_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10991_ _03827_ _03832_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12730_ _05607_ _05608_ _05609_ _05610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_96_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12661_ _05533_ _05534_ _05535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11612_ _04452_ _04453_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12592_ _02499_ _00397_ _05415_ _05459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12602__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11543_ _04293_ _04306_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_53_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_151_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11474_ _04314_ _04315_ _04316_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_13213_ _06047_ _06048_ _06046_ _06132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10425_ _00388_ _06730_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08034__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07694__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13144_ _00369_ _03725_ _06057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07093__I0 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10356_ _03230_ _03234_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12118__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13075_ _05884_ _05894_ _05983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10287_ _03025_ _03084_ _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_100_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12026_ _04116_ _04867_ _04868_ _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07545__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12928_ _05643_ _05824_ _05825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07848__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11644__A3 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12859_ _02762_ _00397_ _05704_ _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_28_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08050_ _00949_ _00950_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10080__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07001_ _05647_ _05485_ _06640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_77_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09222__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11580__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08952_ net95 _06627_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07903_ net91 net142 _06598_ _06618_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09525__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08883_ _01774_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07536__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11332__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07834_ _00730_ _00735_ _00733_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07765_ _00698_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09289__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13085__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09504_ _02391_ _02392_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07696_ _00659_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09435_ _00370_ _06691_ _02249_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_137_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09366_ _02198_ _02201_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11399__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08317_ _01218_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09297_ _06659_ _00385_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10071__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08248_ _00355_ _05833_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08179_ _06179_ _00373_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08016__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10933__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10210_ _03090_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13529__B _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11190_ _04012_ _04032_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_132_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11571__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10141_ _02998_ _02999_ _03021_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07527__B _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10072_ _02608_ _02704_ _02953_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07527__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12520__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13900_ _00231_ net36 clknet_leaf_19_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_98_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13831_ _00162_ clknet_leaf_44_clk DDS_Stage.xPoints_Generator1.RegF\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10974_ _03816_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13762_ _00097_ clknet_leaf_12_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12823__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12713_ _05558_ _05590_ _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13693_ _00028_ clknet_leaf_6_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12644_ _05421_ _05514_ _05515_ _05516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12575_ _05440_ _05277_ _05441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11526_ _04366_ _04367_ _04368_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_81_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11457_ _04297_ _04298_ _04299_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_124_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10408_ _00398_ _06708_ _06710_ _00394_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11388_ net87 _02236_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10339_ _03217_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13127_ _06037_ _06038_ _06040_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13058_ _05889_ _05963_ _05964_ _05965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12009_ _04850_ _04851_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_108_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07550_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[2\] _00546_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12814__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07481_ _05583_ _06754_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09220_ _00355_ _06701_ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12578__A1 _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09151_ _01990_ _02043_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08102_ _00355_ net152 net155 net58 _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09082_ _01881_ _01941_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09994__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08033_ _06179_ _00376_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08954__B1 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09984_ _02865_ _02866_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08935_ _01825_ _01829_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07509__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08866_ _01757_ _01761_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07817_ _00724_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08797_ _05280_ _01693_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07748_ net112 DDS_Stage.xPoints_Generator1.RegP\[-10\] _00684_ _00690_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10816__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07679_ DDS_Stage.xPoints_Generator1.RegFrequency\[-4\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-4\]
+ _00644_ _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_101_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09418_ _02163_ _02223_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10690_ _03498_ _03512_ _03564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09349_ _02165_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13230__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12360_ _05202_ _05203_ _05208_ _05209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_90_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10044__A2 _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11311_ _00354_ _02940_ _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12291_ _04378_ _04383_ _05134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11242_ _04081_ _04084_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_121_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11173_ _03922_ _03928_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10124_ _02860_ _03004_ _03005_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_101_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06971__A2 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10055_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[19\] _02938_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_54_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13049__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13814_ _00145_ net36 clknet_leaf_47_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_3_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10807__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13745_ _00080_ net36 clknet_leaf_52_clk DDS_Stage.xPoints_Generator1.CosNew\[-8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08476__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10957_ _03795_ _03798_ _03799_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13676_ _00011_ clknet_leaf_3_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10888_ _03727_ _03758_ _05171_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12627_ _05493_ _05497_ _05498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_42_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_42_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09976__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12558_ _02938_ _00381_ _05423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11783__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11509_ _04348_ _04351_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12489_ _05326_ _05345_ _05349_ _05350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_1_clk_I clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07167__B _06782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08400__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ _05420_ _05973_ _06623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_119_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13288__A2 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08720_ _01543_ _01544_ _01542_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08651_ _01477_ _01501_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09900__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07911__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07602_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-15\] DDS_Stage.xPoints_Generator1.RegFrequency\[-15\]
+ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08582_ _06308_ _06179_ _00398_ _00394_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_77_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12799__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07533_ _05409_ _05420_ _06092_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_89_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13460__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11471__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ _06232_ _05572_ _05886_ _06624_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_29_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09203_ _02090_ _02094_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_63_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07395_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-25\] _00418_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_29_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone14_I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09134_ _00355_ _06696_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12971__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09065_ _01868_ _01952_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_116_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08016_ _06618_ _00373_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_130_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07792__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09967_ net53 _02757_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08918_ _01729_ _01733_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09898_ _02779_ _02780_ _02781_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_97_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08849_ _00398_ net155 _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07902__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07902__B2 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11860_ _04694_ _04695_ _04696_ _04702_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_58_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10811_ _03681_ _03673_ _03682_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_28_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11791_ _04628_ _04631_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13451__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13530_ _06323_ _06398_ _06401_ _06474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10742_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[2\] _03609_ _03615_ _03616_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_67_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13461_ _06398_ _06399_ _06400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_138_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10673_ _03472_ _03480_ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_82_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12412_ _04861_ _04871_ _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_153_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13392_ _06324_ _06325_ _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12343_ _05167_ _05189_ _05190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_62_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12274_ _05104_ _05116_ _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_65_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11225_ _03806_ _03811_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_121_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08394__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07197__A2 _06759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11156_ _03985_ _03998_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_147_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10107_ _02980_ _02988_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11087_ _03919_ _03929_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10038_ _02919_ _02920_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11989_ _04773_ _04831_ _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11048__A4 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13728_ _00063_ net36 clknet_leaf_37_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_128_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07121__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13659_ _05822_ _06611_ _06612_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11205__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-19\] _06794_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12705__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09821_ _02701_ _02705_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09752_ _00385_ _06685_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06964_ _05409_ _05908_ _06566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08137__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08703_ _01540_ _01600_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06895_ _05280_ _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_20
X_09683_ _02562_ _02569_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08688__A2 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10495__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08634_ _01530_ _01531_ _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08565_ _01383_ _01384_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_25_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07516_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-3\] _00517_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08496_ _00398_ _05864_ _00394_ _06179_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07112__A2 _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07447_ _06795_ _05995_ _06826_ _05658_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_91_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08860__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06871__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07378_ _00409_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09117_ _02005_ _02009_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_98_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09048_ _01881_ _01941_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_60_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10941__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11010_ _03835_ _03845_ _03815_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10183__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08128__A1 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12961_ _02854_ _00397_ _05805_ _05859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08679__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09876__A1 _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11912_ _00390_ _01956_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11683__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12892_ _03340_ _00378_ _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11843_ net70 _01430_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_67_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10238__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11435__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11774_ _04615_ _04616_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_138_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07103__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13513_ _06385_ _06434_ _06455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10725_ _03515_ _03597_ _03598_ _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_138_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13444_ _06379_ _06380_ _06381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10656_ _03449_ _03457_ _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10587_ _03381_ _03461_ _03462_ _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_140_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13375_ _06305_ _06283_ _06306_ _06307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12326_ _00397_ _01249_ _04405_ _05172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07429__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12257_ _05091_ _05099_ _05100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08367__A1 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11208_ _04043_ _04044_ _04050_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12188_ _05030_ _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_11139_ _03932_ _03945_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08119__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13663__A2 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11269__A4 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_82_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08350_ _00874_ _00875_ _01250_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_86_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07301_ _00353_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11977__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08281_ _00933_ _00937_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_18_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13179__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07232_ _05182_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-10\] _00297_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_4_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ _05409_ _06651_ _05875_ _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_70_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10401__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07948__A4 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07094_ _06719_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06908__A2 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ _02612_ _02620_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11901__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07030__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ _00897_ _00893_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_66_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09735_ _02595_ _02612_ _02620_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06947_ _05778_ _06373_ _06383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08125__A4 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09666_ _02460_ _02551_ _02552_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06878_ _05627_ _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_124_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08617_ _01213_ _01238_ _01335_ _01336_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA__13894__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12209__A3 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09597_ _02479_ _02483_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_3_4__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11417__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08548_ _01445_ _01446_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11968__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07097__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08479_ _01264_ _01265_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_65_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10510_ _03302_ _03385_ _03386_ _03387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11490_ _04330_ _04331_ _04332_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_80_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12917__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10441_ _03138_ _03226_ _03225_ _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09389__A3 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08597__B2 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13160_ _06069_ _06074_ _06075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10372_ _03107_ _03165_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12111_ _00397_ _01610_ _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13091_ _05981_ _05985_ _06000_ _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_130_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12042_ _04882_ _04883_ _04884_ _04885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12944_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-9\] _05841_ _05842_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_clkbuf_leaf_56_clk_I clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13885__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12875_ _05764_ _05765_ _05766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07875__A3 _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11826_ _04666_ _04667_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07088__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11757_ _04538_ _04598_ _04599_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_155_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10708_ _03581_ _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_155_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11688_ _00372_ _01249_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12908__A1 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13427_ _06302_ _06363_ _06364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10639_ _03452_ _03455_ _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08588__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12384__A2 _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08588__B2 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13358_ _06288_ _06289_ _06290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_122_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12309_ _05147_ _05152_ net65 _05153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07260__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13289_ _06212_ _06213_ _06214_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12687__A3 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07012__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10698__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ _06179_ _00379_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11895__A1 _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07175__B _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08760__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08760__B2 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07781_ _00706_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13636__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 net109 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09520_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[13\] _02409_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_127_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11647__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08512__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13876__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09451_ _02291_ _02299_ _02339_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_149_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08402_ _00909_ _00924_ _01302_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_149_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09382_ _02263_ _02271_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_148_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_35_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08333_ _01234_ _01199_ _01211_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XPHY_EDGE_ROW_49_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12611__A3 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10083__B1 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08264_ _01096_ _01144_ _01165_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07215_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-13\] _06822_ _06823_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08195_ _05864_ _00370_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08579__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ _06764_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10386__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13800__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07077_ _05409_ _06651_ _06704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_58_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10138__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07085__B _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08751__A1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07979_ _00857_ _00860_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09718_ _02601_ _02602_ _02603_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10990_ _03827_ _03832_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_97_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08503__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13867__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09649_ _02534_ _02535_ _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10310__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12660_ _05438_ _05445_ _05534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_104_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11611_ _04452_ _04453_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_136_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12591_ _05456_ _05457_ _05458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11542_ _04375_ _04384_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_136_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07490__A1 _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11473_ _00378_ _01792_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13212_ _05740_ _06034_ _06127_ _06130_ _06131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_150_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10424_ _00382_ _06742_ _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_150_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13143_ _05958_ _05959_ _05953_ _06056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10355_ _03231_ _03232_ _03233_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_EDGE_ROW_76_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13315__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12118__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13074_ _05888_ _05982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10286_ _03107_ _03165_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12025_ _04117_ _04118_ _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11877__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08742__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07545__A2 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13858__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12927_ _05719_ _05824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_85_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11644__A4 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12858_ _05701_ _05703_ _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_28_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11809_ _00372_ _01247_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12789_ _05670_ _05671_ _05672_ _05673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_32_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07481__A1 _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07000_ _05409_ _05572_ _06639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_94_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09222__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10368__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07233__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08951_ _00352_ _06691_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07902_ net91 _06598_ _06618_ net143 _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08882_ _01513_ _01518_ _01777_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11332__A3 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09930__B1 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07833_ _00733_ _00734_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10540__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07764_ net6 DDS_Stage.xPoints_Generator1.RegP\[-2\] _00684_ _00698_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09289__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09503_ _02320_ _02321_ _02390_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__13849__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07695_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-2\] _00658_ _00395_ _00659_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clone44_I net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ _02322_ _02248_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12045__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09365_ _02182_ _02190_ _02254_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08316_ _01216_ _01204_ _01217_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09296_ _06654_ _00388_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08247_ net73 _05398_ _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07472__A1 _06799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07472__B2 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08178_ _01078_ _01079_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07224__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _05897_ _06748_ _06749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10140_ _03020_ _02997_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10071_ net95 _06696_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12520__A2 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13830_ _00161_ clknet_leaf_45_clk DDS_Stage.xPoints_Generator1.RegF\[-3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13761_ _00096_ clknet_leaf_78_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10973_ _00378_ net135 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12712_ _05576_ _05589_ _05590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13692_ _00027_ clknet_leaf_8_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12643_ _05422_ _05423_ _05515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_155_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12574_ _04036_ _04104_ _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11525_ _00361_ _02238_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11456_ _00359_ _02238_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07215__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10407_ _02704_ _03283_ _03284_ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11387_ net83 _02153_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13126_ _05280_ net33 _06040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10338_ _03142_ _03150_ _03216_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10770__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13057_ _05890_ _05891_ _05964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10269_ _03146_ _03147_ _03148_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_84_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12008_ _04115_ _04119_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07480_ _00488_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09150_ _01992_ _02042_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10589__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08101_ _00992_ _01001_ _01002_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07454__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09081_ _01969_ _01973_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08032_ _06308_ _00373_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07206__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08954__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08954__B2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ _02787_ _02795_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08934_ _01826_ _01827_ _01828_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07509__A2 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08865_ _01758_ _01759_ _01760_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10513__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07816_ _00382_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[25\] _00395_ _00724_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08796_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[5\] _01693_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07747_ _00689_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_154_Right_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07678_ _00642_ _00643_ _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_101_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09417_ _02163_ _02223_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09348_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[12\] _02238_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_118_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09279_ _02168_ _02169_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_105_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11310_ _00351_ _03018_ _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12290_ _04401_ _04406_ _05132_ _05133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11241_ _04082_ _04083_ _03855_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_132_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08945__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11172_ _03960_ _03965_ _04014_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_30_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10123_ _02863_ _02922_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10054_ _05182_ _02936_ _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09370__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13813_ _00144_ net36 clknet_leaf_50_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_3_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10807__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13744_ _00079_ net36 clknet_leaf_67_clk DDS_Stage.xPoints_Generator1.CosNew\[-9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_74_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10956_ _03796_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_86_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13675_ _00010_ clknet_leaf_77_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10887_ _03729_ _03754_ _03757_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_128_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12626_ _05494_ _05495_ _05497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07436__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12557_ _02854_ _00384_ _05422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11508_ _04350_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12488_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-15\] _05281_ _05348_ _05349_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11439_ _04276_ _04281_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_110_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13109_ _05250_ _06016_ _06018_ _06020_ _06021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_06980_ _05409_ _06621_ _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_95_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08650_ _01546_ _01547_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07183__B _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07601_ _00577_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07911__A2 _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08581_ _06179_ _00398_ _00394_ _06308_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09113__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12799__A2 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07532_ _00530_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07463_ _06778_ _06787_ _05658_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11471__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09202_ _02091_ _02092_ _02093_ _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_92_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ _00417_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07427__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09133_ _01927_ _01935_ _02025_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_20_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12971__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ _06059_ _01955_ _01957_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_116_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10982__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08015_ _00912_ _00916_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11931__B1 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09966_ _02848_ _02849_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_08917_ _01737_ _01766_ _01811_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09897_ net60 _06742_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08848_ _01667_ _01742_ _01743_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07902__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08779_ net60 _06664_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10939__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10810_ _03668_ _03669_ _03667_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_28_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11790_ _04617_ _04618_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_68_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10741_ _03612_ _03614_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13460_ _00378_ _03727_ _06324_ _06399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10672_ _03546_ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_137_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12411_ _05262_ _05263_ _05264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07418__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13391_ _00378_ _03725_ _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone31 net136 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_91_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone53 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-20\] net152 vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlya_4
Xclkbuf_leaf_20_clk clknet_3_6__leaf_clk clknet_leaf_20_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12342_ _05176_ _05187_ _05188_ _05189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08091__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12273_ _05108_ _05115_ _05116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11224_ _04057_ _04065_ _04066_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08394__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11155_ _03997_ _03993_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_147_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10106_ _02983_ _02987_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11086_ _03922_ _03928_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10037_ _00370_ _06738_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11988_ _04772_ _04775_ _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13727_ _00062_ net36 clknet_3_3__leaf_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10939_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-2\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-2\]
+ _05171_ _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13658_ _05280_ net26 _06612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12609_ _05472_ _05477_ _05478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07409__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11205__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13589_ _06535_ _06536_ _06537_ _06538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xclkbuf_leaf_11_clk clknet_3_6__leaf_clk clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10964__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12705__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09820_ _02608_ _02702_ _02704_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_111_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09751_ _00388_ _06679_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06963_ _05572_ _06092_ _06555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_78_clk clknet_3_2__leaf_clk clknet_leaf_78_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08137__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08702_ _01548_ _01550_ _01599_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_09682_ _02567_ _02568_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06894_ _05387_ _05756_ _05800_ _05811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08633_ _01422_ _01424_ _01437_ _01506_ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08564_ _01459_ _01462_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_25_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07515_ _00516_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08495_ _01287_ _01393_ _01394_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_49_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout36 net19 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_0_76_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07446_ _06713_ _05897_ _06070_ _06721_ _05658_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08860__A3 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07377_ DDS_Stage.xPoints_Generator1.CosNew\[-9\] DDS_Stage.xPoints_Generator1.RegP\[-9\]
+ _00402_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06871__A2 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09116_ _02006_ _02007_ _02008_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_98_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07820__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09047_ _01889_ _01940_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09573__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10183__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_129_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09949_ _02769_ _02832_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10242__B net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_69_clk clknet_3_0__leaf_clk clknet_leaf_69_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08128__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12960_ _05803_ _05804_ _05858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11911_ _00397_ _01792_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_142_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12891_ _05670_ _05782_ _05783_ _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12880__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11683__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11842_ net54 _01524_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_clk_I clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11435__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11773_ _00361_ _01524_ _01430_ _00365_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07270__C _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13512_ _06453_ _06446_ _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10724_ _03518_ _03526_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_95_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13443_ _06229_ _06360_ _06380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10655_ _03449_ _03457_ _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_64_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13374_ _06234_ _06282_ _06306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10586_ _03384_ _03393_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10946__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12325_ _04391_ _05168_ _05169_ _05170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12148__B1 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12256_ _05093_ _05098_ _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08367__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11207_ _04045_ _04049_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09564__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13360__A2 _06208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12187_ _05027_ _05028_ _05029_ _05030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_76_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11138_ _03948_ _03967_ _03980_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08119__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11069_ _03896_ _03898_ _03911_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
Xclkbuf_leaf_0_clk clknet_3_2__leaf_clk clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_69_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07878__A1 _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12623__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07300_ net66 net58 _05182_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08280_ _01077_ _01082_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_6_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13179__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07231_ _05658_ _06125_ _06749_ _00295_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_61_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07162_ _05409_ _05789_ _06778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07802__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07093_ _06710_ _06718_ _05182_ _06719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09555__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09803_ _02620_ _02612_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__07030__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ _00894_ _00895_ _00896_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XPHY_EDGE_ROW_105_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09734_ _02535_ _02619_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06946_ _05420_ _05496_ _05409_ _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__11114__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07869__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09665_ _02461_ _02462_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06877_ _05387_ _05398_ _05616_ _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ _01233_ _01235_ _01213_ _01514_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_94_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09596_ _02479_ _02483_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__12209__A4 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11417__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08547_ _06633_ _00373_ _01377_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07798__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07097__A2 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08478_ _01374_ _01377_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07429_ _05886_ _06754_ _06646_ _05658_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_114_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12917__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10440_ _03218_ _03316_ _03317_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__A4 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08597__A2 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10371_ _03110_ _03164_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12110_ _04949_ _04952_ _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13090_ _05990_ _05999_ _06000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09546__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12041_ _00393_ _01792_ _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11353__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_123_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12943_ _05829_ _05840_ _05841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12874_ net86 net54 _03727_ _05765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_87_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07875__A4 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11825_ _04666_ _04667_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12605__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11756_ _04586_ _04597_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_138_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10707_ _03577_ _03580_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11687_ _04526_ _04529_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13426_ _06304_ _06361_ _06363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12908__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10638_ _03498_ _03512_ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13030__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10919__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08588__A2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13357_ _06217_ _06218_ _06286_ _06289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_10569_ _03387_ _03444_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12308_ _04371_ _04385_ _05152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13288_ _05280_ net35 _06214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09537__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12239_ _05079_ _05080_ _05081_ _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_20_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12687__A4 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07012__A2 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10698__A3 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08760__A2 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07780_ DDS_Stage.xPoints_Generator1.RegFrequency\[-9\] DDS_Stage.xPoints_Generator1.RegF\[-9\]
+ _00402_ _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput4 net127 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11647__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12844__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08512__A2 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09450_ _02277_ _02290_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_149_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08401_ _00394_ _05398_ _00844_ _00923_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09381_ _02266_ _02270_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08332_ _01175_ _01176_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07323__I0 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12611__A4 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10083__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10083__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08263_ _01121_ _01142_ _01164_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07214_ _06819_ _06820_ _06821_ _05658_ _05171_ _06822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_85_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08194_ _01095_ _00983_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_43_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08579__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07145_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-24\] _06758_ _06763_
+ _06764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_131_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11583__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07076_ _05572_ _05452_ _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_112_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10138__A2 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11335__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08200__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08751__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07554__A3 _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ _00846_ _00863_ _00879_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09717_ _00363_ _06730_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06929_ _05822_ _06179_ _06190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08503__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09648_ _06664_ _06659_ _00398_ _00394_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__10310__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09579_ _02448_ _02466_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_104_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11610_ _04234_ _04235_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_46_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12590_ _05408_ _05427_ _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07314__I0 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11541_ _04378_ _04383_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13012__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11472_ _00372_ _01956_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13211_ _06122_ _06128_ _06129_ _06033_ _06119_ _06130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_122_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10423_ _03231_ _03299_ _03300_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11574__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10377__A2 _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13142_ _06053_ _06054_ _06055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10354_ _00385_ _06730_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09519__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13315__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13073_ _05910_ _05918_ _05980_ _05981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10285_ _03110_ _03164_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12024_ _04117_ _04118_ _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11877__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08742__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13079__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12926_ _05741_ _05821_ _05823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12857_ _05695_ _05744_ _05746_ _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11808_ _00372_ _01247_ _04650_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_12788_ _00361_ _03558_ _05672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11739_ _04577_ _04581_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13003__A1 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07481__A2 _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13409_ _06275_ _06277_ _06344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_25_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07233__A2 _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13794__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08950_ _00355_ _06685_ _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07901_ _00789_ _00797_ _00802_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08881_ _01425_ _01507_ _01605_ _01687_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07832_ _00731_ _00732_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09930__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11332__A4 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09930__B2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10540__A2 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07763_ _00697_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09502_ _02320_ _02321_ _02390_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08497__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07694_ DDS_Stage.xPoints_Generator1.CosNew\[-2\] _00657_ _00577_ _00658_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09433_ _02246_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09364_ _02185_ _02189_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13242__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12045__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08315_ _01182_ _01183_ _01203_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10056__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09295_ _06664_ _00382_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08246_ _01127_ _01130_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_105_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08177_ _05833_ _00379_ _00376_ _05864_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11556__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_55_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07128_ _05572_ _05431_ _05409_ _06748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__07224__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13785__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07096__B _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07059_ _06687_ _06688_ _06689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11308__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10070_ _02876_ _02878_ _02951_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09921__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13760_ _00095_ clknet_leaf_78_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10972_ _03806_ _03811_ _03814_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10295__A1 _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12711_ _05579_ _05588_ _05589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13691_ _00026_ clknet_leaf_8_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12642_ _05422_ _05423_ _05514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10047__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09988__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12573_ _04105_ _04174_ _05439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_80_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__B1 _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11524_ _00365_ _02236_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07463__A2 _06787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08660__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11455_ _00351_ _02499_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10406_ net63 _06710_ net57 _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11386_ _04226_ _04227_ _04228_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13125_ _06029_ _06033_ _06035_ _05182_ _06038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_10337_ _03145_ _03215_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06974__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10770__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13056_ _05890_ _05891_ _05963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_72_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10268_ _00385_ _06724_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12007_ _04832_ _04837_ _04849_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10199_ _03078_ _03079_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13472__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12909_ _02940_ _00390_ _05804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07151__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13889_ _00220_ net36 clknet_leaf_9_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_33_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08100_ _00996_ _01000_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11786__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09080_ _01970_ _01971_ _01947_ _01972_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_71_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08031_ _00757_ _00932_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11538__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07206__A2 _06811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08954__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09982_ _02775_ _02786_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06965__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06965__B2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08933_ _06637_ _00385_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08864_ net60 _06672_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10513__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07815_ _00723_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08795_ _01688_ _01691_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07746_ net118 DDS_Stage.xPoints_Generator1.RegP\[-11\] _00684_ _00689_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07677_ DDS_Stage.xPoints_Generator1.RegFrequency\[-5\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-5\]
+ _00638_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07142__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09416_ _02241_ _02305_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_137_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09347_ _02233_ _02235_ _02237_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09278_ _00370_ _06685_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08229_ _01127_ _01130_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11240_ _00354_ _03018_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08945__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11171_ _03955_ _04013_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10122_ _02863_ _02922_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_54_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10053_ _02929_ _02934_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10504__A2 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09370__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13930__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13812_ _00143_ net36 clknet_leaf_50_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_3_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10268__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13743_ _00078_ net36 clknet_leaf_68_clk DDS_Stage.xPoints_Generator1.CosNew\[-10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10955_ _03796_ _03797_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07133__A1 _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13206__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10886_ _03677_ _03721_ _03755_ _03756_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13674_ _00009_ clknet_leaf_1_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12625_ _03266_ _00372_ _05495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07436__A2 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12556_ _02762_ _00387_ _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11507_ _04336_ _04337_ _04349_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12487_ _05339_ _05347_ _05340_ _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_80_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11438_ _04277_ _04278_ _04280_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_123_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10155__B _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13749__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11369_ _04181_ _04182_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06947__A1 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11940__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13108_ _05629_ _05831_ _06019_ _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_13039_ _02938_ _00397_ _05909_ _05944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07464__B _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13921__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07600_ DDS_Stage.LCU.SelMuxConfigReg _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08580_ _01402_ _01404_ _01478_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10259__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09113__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07531_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-1\] _00529_ _00530_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07124__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07462_ _05897_ _06666_ _05409_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09201_ _06654_ _00385_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07393_ DDS_Stage.xPoints_Generator1.CosNew\[-1\] DDS_Stage.xPoints_Generator1.RegP\[-1\]
+ _00402_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09132_ _01930_ _01934_ _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09063_ _05280_ _01956_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08014_ _00913_ _00914_ _00915_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10982__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12184__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06938__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11931__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11931__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09965_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-8\] _02847_ _02849_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08916_ _01740_ _01765_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09896_ net61 _06738_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08847_ _01668_ _01669_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13912__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ net91 _06659_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13436__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07729_ _00679_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10740_ _03476_ _03479_ _03613_ _03472_ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__08863__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10670__B2 _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ _03413_ _03481_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12410_ _05254_ _05255_ _05263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclone10 net88 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13390_ _06322_ _06323_ _06324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_129_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclone21 net78 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xclone43 net144 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_12341_ _05185_ _05186_ _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclone54 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-20\] net153 vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlya_4
XFILLER_0_145_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08091__A2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__A2 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12272_ _05110_ _05114_ _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_121_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11223_ _04063_ _04064_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06929__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11154_ _03994_ _03995_ _03996_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_8_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10105_ _02984_ _02985_ _02986_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_65_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11085_ _03924_ _03927_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10489__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10036_ _02916_ _02918_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13903__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11987_ _04803_ _04828_ _04829_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13726_ _00061_ net36 clknet_leaf_24_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_129_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10938_ _03785_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10869_ _03696_ _03714_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13657_ _06606_ _06610_ _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_128_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12608_ _05473_ _05475_ _05476_ _05477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__07409__A2 _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13588_ _00390_ _03679_ _06537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12539_ _05399_ _05400_ _05401_ _05402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_26_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10964__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09031__A1 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11913__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07593__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06962_ _06059_ _06513_ _06534_ _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09750_ _00382_ _06691_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08701_ _01571_ _01598_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09681_ _00370_ _06708_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06893_ _05767_ _05778_ _05789_ _05800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08632_ _01437_ _01506_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08563_ _01460_ _01461_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07514_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-4\] _00515_ _00395_ _00516_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_25_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08494_ _01288_ _01289_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_76_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07445_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-16\] _00459_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_135_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08860__A4 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07376_ _00408_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09115_ _06649_ _00385_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11601__B1 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09046_ _01891_ _01939_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07820__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09573__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09948_ _02822_ _02831_ _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_129_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09879_ _02760_ _02761_ _02763_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11910_ _04747_ _04752_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_142_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12890_ _05671_ _05672_ _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12880__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11841_ net66 _01610_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11772_ _00361_ _00365_ _01524_ _01430_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__08836__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10723_ _03518_ _03526_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_27_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13511_ _06381_ _06436_ _06453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10654_ _03496_ _03528_ _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_126_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13442_ _06307_ _06359_ _06379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13373_ _06231_ _06305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10585_ _03384_ _03393_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_50_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12324_ _04393_ _04407_ _05169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_51_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12148__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12148__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12255_ _05096_ _05097_ _05098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09013__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11206_ _04046_ _04047_ _04048_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_103_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09564__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12186_ _00390_ _01610_ _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XDDS_Module_50 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_11137_ _03918_ _03947_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11068_ _03902_ _03910_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_69_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10019_ _02813_ _02901_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07878__A2 _06523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08827__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12623__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10634__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13709_ _00044_ clknet_leaf_33_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07230_ _05409_ _00294_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06872__I _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12387__A1 _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-21\] _06777_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_15_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07092_ _05658_ _06717_ _06718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09004__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09555__A2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09802_ _02685_ _02686_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07994_ _00363_ _06637_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06945_ _05409_ _06351_ _06362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09733_ _02615_ _02618_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11114__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07869__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06876_ _05171_ _05540_ _05605_ _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09664_ _02461_ _02462_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10873__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08615_ _01096_ _01144_ _01238_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_124_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09595_ _02325_ _02481_ _02482_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_124_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12075__B1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08546_ _01375_ _01376_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_77_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10625__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08477_ _01375_ _01376_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_147_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09491__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ _06059_ _00440_ _00445_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07359_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-1\] _00398_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_0_73_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_149_Right_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10370_ _03191_ _03194_ _03248_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_131_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09029_ _01848_ _01856_ _01922_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_130_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12040_ _00390_ _01794_ _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07319__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09546__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07557__A1 _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07546__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11353__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12550__A1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07309__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12942_ _05336_ _05834_ _05835_ _05839_ _05840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12873_ net66 net54 _03727_ _05764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11824_ _04632_ _04633_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12605__A2 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10616__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11755_ _04586_ _04597_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09482__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10706_ _03037_ _03579_ _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07493__B1 _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11686_ _04527_ _04528_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13425_ _06229_ _06360_ _06361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10637_ _03505_ _03511_ _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07245__B1 _06732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10568_ _03391_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13356_ _06217_ _06218_ _06286_ _06288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_52_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12307_ _05133_ _05135_ _05136_ _05151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_87_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10499_ _03287_ _03375_ _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13287_ _06131_ _06210_ _05182_ _06213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09537__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12238_ _00361_ _02409_ _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07548__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12169_ _04934_ _04935_ _04913_ _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__10698__A4 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 net132 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10855__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08400_ _06633_ _00370_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09380_ _02267_ _02268_ _02269_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_148_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08331_ _01171_ _01231_ _01232_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_35_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07323__I1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10083__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08262_ _01139_ _01141_ _01145_ _01163_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11280__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07213_ _06713_ _06681_ _06748_ _05496_ _06821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_08193_ _01069_ _01094_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__09225__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07144_ _06760_ _06762_ _05171_ _06763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_95_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11032__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08579__A3 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11583__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07075_ _06059_ _06700_ _06702_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11335__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08200__A2 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07977_ _00848_ _00862_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09716_ _00367_ _06724_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11099__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06928_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-22\] _06179_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08503__A3 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09647_ _06659_ _00398_ _00394_ _06664_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06859_ DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[0\] _05431_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_97_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09578_ _02451_ _02465_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_104_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08529_ _05182_ _01428_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_46_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09464__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07314__I1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11540_ _04379_ _04380_ _04382_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07475__B1 _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11471_ _00375_ _01794_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_137_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13012__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10422_ _03232_ _03233_ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13210_ _06030_ _06119_ _06120_ _06129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_21_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11574__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10353_ _00388_ _06724_ _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13141_ _05961_ _05976_ _06054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_150_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13072_ _05913_ _05979_ _05980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _03154_ _03163_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12023_ _04848_ _04852_ _04865_ _04866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__13079__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07950__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12925_ _05743_ _05820_ _05821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_87_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12856_ _05699_ _05715_ _05746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_38_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11807_ _04646_ _04649_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_84_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09455__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12787_ _03556_ _00365_ _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11738_ _04579_ _04580_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_154_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13003__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11669_ _04460_ _04461_ _04440_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_98_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11014__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13408_ _06275_ _06277_ _06343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07218__B1 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13339_ _06268_ _06269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_51_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_90_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07900_ _00792_ _00796_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08880_ _01699_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07831_ _00731_ _00732_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09930__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07941__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07762_ net5 DDS_Stage.xPoints_Generator1.RegP\[-3\] _00684_ _00697_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09501_ _02325_ _02327_ _02389_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_116_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_142_Left_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07693_ DDS_Stage.xPoints_Generator1.RegFrequency\[-2\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-2\]
+ _00656_ _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08497__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09432_ _02241_ _02305_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09363_ _02192_ _02220_ _02252_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13242__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12045__A3 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08314_ _01182_ _01183_ _01203_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10056__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09294_ _02091_ _02183_ _02184_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08245_ _01124_ _01132_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08176_ _05864_ _05833_ _00379_ _00376_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_31_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11556__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07127_ _05658_ _05540_ _06746_ _06747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07224__A3 _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07058_ _05409_ _06125_ _06688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_2_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11308__A2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06983__A2 _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09921__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10971_ _03813_ _03805_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12710_ _05581_ _05587_ _05588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11492__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13690_ _00025_ clknet_leaf_10_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07160__A2 _06776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12641_ _05509_ _05512_ _05513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10047__A2 _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09988__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12572_ _05434_ _05437_ _05438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__07999__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07999__B2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11523_ _00369_ _02153_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08660__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11454_ _00354_ _02409_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10405_ net63 _06710_ net57 _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11385_ net66 net54 _02153_ _02051_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_59_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07287__B _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13124_ _06030_ _06036_ _06037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10336_ _03149_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13055_ _05954_ _05960_ _05961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10267_ _00388_ _06710_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_72_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08176__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12006_ _04835_ _04836_ _04849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10198_ _03073_ _03074_ _03077_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07923__A1 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13957_ _00288_ net36 clknet_leaf_58_clk DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__13472__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12908_ _02938_ _00393_ _05803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13888_ _00219_ net36 clknet_leaf_37_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07151__A2 _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12839_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-11\] _05631_ _05728_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11235__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11786__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08030_ _00931_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_154_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06880__I _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11538__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09981_ _02799_ _02820_ _02797_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_122_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06965__A2 _06081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08932_ _06633_ _00388_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08863_ net92 _06664_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_150_Left_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07814_ _00379_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[24\] _00395_ _00723_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08794_ _01529_ _01689_ _01690_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07745_ _00688_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13662__B _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09667__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07676_ DDS_Stage.xPoints_Generator1.RegFrequency\[-5\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-5\]
+ _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07142__A2 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09415_ _02243_ _02304_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_101_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09346_ _05280_ _02236_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09277_ _02165_ _02167_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_134_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08228_ _01102_ _01129_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08159_ _01060_ _01057_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_28_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11170_ _03959_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08945__A3 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10121_ _02943_ _03002_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_98_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07327__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10052_ _02929_ _02934_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07905__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13811_ _00142_ net36 clknet_leaf_52_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_145_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10268__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13742_ _00077_ net36 clknet_leaf_68_clk DDS_Stage.xPoints_Generator1.CosNew\[-11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10954_ _00381_ _02499_ _02409_ _00384_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_85_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13673_ _00008_ clknet_leaf_0_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10885_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[4\] _03720_ _03756_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11217__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12624_ _03189_ _00375_ _05494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06892__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12555_ _04026_ _05417_ _05418_ _05419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10976__B1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11506_ _00397_ _01247_ _04338_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_145_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12486_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-17\] _05341_ _05347_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11437_ _04279_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11368_ _04175_ _04210_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06947__A2 _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11940__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13107_ _05725_ _05836_ _05838_ _06019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10319_ _03121_ _03129_ _03197_ _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08149__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11299_ _04047_ _04048_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_119_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13038_ _05906_ _05907_ _05943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09897__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11456__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07530_ _05171_ _00527_ _00528_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_89_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10259__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_54_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07124__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07461_ _00471_ _00472_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09200_ _06649_ _00388_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06883__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07392_ _00416_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09131_ _01918_ _02023_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08085__B1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_69_clk_I clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09062_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[8\] _01956_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_114_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08013_ _06308_ _00385_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08388__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12184__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11931__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07060__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09964_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-8\] _02847_ _02848_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08915_ _01808_ _01809_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09895_ net73 _06744_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11695__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ _01668_ _01669_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08560__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08777_ net73 _06672_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07728_ net4 DDS_Stage.xPoints_Generator1.RegF\[-4\] _00667_ _00679_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07659_ DDS_Stage.xPoints_Generator1.CosNew\[-7\] _00627_ _00577_ _00628_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08863__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10670_ _03345_ net79 _03343_ _02681_ _03350_ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_36_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12947__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09329_ _02194_ _02219_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclone11 net64 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_152_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09812__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclone22 net146 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_129_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone44 net144 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_106_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12340_ _05185_ _05186_ _05187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12271_ _05112_ _05113_ _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08379__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11222_ _04063_ _04064_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_120_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06929__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07051__A1 _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11153_ _00365_ _03266_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_147_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10104_ _00385_ _06708_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11084_ _03925_ _03926_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10035_ _02805_ _02806_ _02917_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10489__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11986_ _04815_ _04827_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13725_ _00060_ net36 clknet_leaf_16_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_TAPCELL_ROW_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10937_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-3\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-3\]
+ _05171_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06865__A1 _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13656_ _06511_ _06607_ _06608_ _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10868_ _03699_ _03713_ _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12607_ net66 _03679_ _05476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13587_ _00393_ _03558_ _06536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10799_ _03612_ _03614_ _03609_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12538_ _03189_ _00372_ _05401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07459__C _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12469_ _04943_ _05016_ _05328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10177__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09031__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11913__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07042__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06961_ _05822_ net155 _06534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08700_ _01574_ _01597_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09680_ _02564_ _02566_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06892_ _05420_ _05485_ _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_55_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08631_ _01435_ _01521_ _01528_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_77_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ _06633_ _00376_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_25_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07513_ _05658_ _00513_ _00514_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08493_ _01288_ _01289_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07444_ _06059_ _00457_ _00458_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07375_ DDS_Stage.xPoints_Generator1.CosNew\[-10\] DDS_Stage.xPoints_Generator1.RegP\[-10\]
+ _00402_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_146_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone12_I net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09114_ _06642_ _00388_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11601__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11601__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07281__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09045_ _01911_ _01938_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07033__A1 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09947_ _02829_ _02830_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_129_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09878_ _05280_ _02762_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09730__B1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08829_ _01723_ _01724_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13897__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11840_ _04680_ _04681_ _04682_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11771_ _04570_ _04583_ _04540_ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08836__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13510_ _06369_ _06443_ _06445_ _06131_ _06451_ _06452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_10722_ _03565_ _03595_ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13441_ _06375_ _06377_ _06378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10653_ _03513_ _03527_ _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_119_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13372_ _06223_ _06284_ _06303_ _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10584_ _03424_ _03459_ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12323_ _04393_ _04407_ _05168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_133_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13345__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12148__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12254_ _04961_ _04963_ _05097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_121_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10159__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09013__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11205_ _00393_ _02153_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07024__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12185_ _00393_ _01524_ _05028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08772__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDDS_Module_40 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XDDS_Module_51 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_11136_ _03977_ _03978_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11067_ _03905_ _03909_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_69_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13888__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10018_ _02812_ _02813_ _02814_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_58_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_82_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11969_ _04809_ _04810_ _04811_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__08827__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13708_ _00043_ clknet_leaf_33_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10634__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13639_ _06586_ _06588_ _06590_ _06591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_116_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07160_ _06771_ _06776_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12387__A2 _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07263__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13812__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07091_ _06712_ _06716_ _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13336__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09004__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10624__B net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07015__A1 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09555__A3 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08763__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09801_ _02644_ _02652_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07810__I0 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10570__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07993_ net74 _06633_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09732_ _02616_ _02617_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06944_ _05583_ _06340_ _06351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09712__B1 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13879__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09663_ _02546_ _02549_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10322__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06875_ _05409_ _05594_ _05605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07869__A3 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08614_ _01326_ _01313_ _01511_ _01243_ _01512_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_124_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09594_ _02480_ _02389_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_124_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08545_ _01369_ _01388_ _01443_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12075__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12075__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10625__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08476_ _06627_ _00376_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09491__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07427_ _06146_ _00442_ _00443_ _00444_ _05280_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_107_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07358_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-1\] _00397_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_0_45_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13803__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07254__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ _00342_ _00343_ _05182_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09028_ _01851_ _01855_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12550__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10561__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07335__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07309__A2 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12941_ _05725_ _05836_ _05837_ _05838_ _05839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XPHY_EDGE_ROW_37_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07562__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12872_ _05762_ _05763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11823_ _04656_ _04664_ _04665_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_64_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11754_ _04592_ _04596_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09482__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10705_ net57 _02704_ _03578_ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_83_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11685_ _00375_ _01249_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08690__B1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13566__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13424_ _06307_ _06359_ _06360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10636_ _03507_ _03510_ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_37_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07245__A1 _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07245__B2 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13355_ _06141_ _06285_ _06286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10567_ _03426_ _03442_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13318__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12306_ _05148_ _05149_ _05150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_23_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13286_ _06131_ _06210_ _06212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_122_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10498_ _03371_ _03374_ _03375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12237_ _00365_ _02238_ _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09537__A3 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10001__B1 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12168_ _04986_ _05009_ _05010_ _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10552__A1 _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11119_ _00393_ _02409_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12099_ _04912_ _04940_ _04941_ _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xinput6 net123 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08330_ _01173_ _01192_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11804__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08261_ _01146_ _01154_ _01161_ _01162_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07484__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11280__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07212_ _05658_ _06755_ _06820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_145_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08192_ _01074_ _01093_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__09225__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07236__A1 _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07143_ _05658_ _06761_ _06762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_95_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11032__A2 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08579__A4 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07074_ _05822_ _06701_ _06702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10791__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11335__A3 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10543__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08200__A3 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07976_ _00840_ _00865_ _00877_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09715_ _00357_ _06738_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06927_ _06114_ _06135_ _06157_ _06168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11099__A2 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _02432_ _02531_ _02532_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10846__A2 _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06858_ DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[2\] _05420_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_20
XANTENNA__08503__A4 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09577_ _02456_ _02464_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08528_ _01320_ _01426_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_104_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09464__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07475__A1 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08459_ _06627_ _00373_ _01270_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07475__B2 _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13548__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13620__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11470_ _04265_ _04311_ _04312_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _03232_ _03233_ _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_61_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07227__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13140_ _05954_ _05960_ _06053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10352_ _00382_ _06738_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13071_ _05917_ _05979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_130_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10283_ _03082_ _03162_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12022_ _04850_ _04851_ _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07950__A2 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12924_ _05751_ _05819_ _05820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_69_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12039__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12855_ _05699_ _05715_ _05744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_38_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11806_ _04647_ _04646_ _04648_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_84_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12786_ _03485_ _00369_ _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09455__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11737_ _04468_ _04470_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_54_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07466__B2 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13539__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11668_ _04509_ _04510_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13407_ _06341_ _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07218__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10619_ _03492_ _03493_ _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07218__B2 _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11014__A2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11599_ _04426_ _04427_ _04428_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13338_ _06263_ _06267_ _06268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13269_ _06174_ _06177_ _06193_ _06194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09391__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07830_ net152 _00376_ _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07941__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07761_ _00696_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09143__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09500_ _02335_ _02388_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_155_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07692_ _00654_ _00655_ _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08497__A3 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09431_ _02243_ _02304_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_121_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_149_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09362_ _02194_ _02219_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12045__A4 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08313_ _00945_ _00978_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__07457__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09293_ _02092_ _02093_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_7_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08244_ _01133_ _01135_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08175_ _05398_ _00382_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_119_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08957__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ _05409_ _05778_ _05789_ _06746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10764__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07057_ _06232_ _06620_ _06687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11308__A3 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10516__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07959_ _00857_ _00860_ _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09134__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10970_ _03796_ _03812_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09629_ _02431_ _02435_ _02515_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11492__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12640_ _05510_ _05511_ _05512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07448__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12441__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-23\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12571_ _03850_ _05435_ _05436_ _05437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09988__A3 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_50_clk clknet_3_1__leaf_clk clknet_leaf_50_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__A2 _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11522_ _04364_ _04360_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_151_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11453_ _04262_ _04294_ _04295_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10404_ _03278_ _03281_ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_34_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11384_ net66 _02153_ _02051_ net54 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10755__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13123_ _06033_ _06035_ _06036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10335_ _03198_ _03213_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07620__A1 DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13054_ _05958_ _05959_ _05960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10266_ _00382_ _06730_ _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08176__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12005_ _04782_ _04785_ _04847_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10197_ _03073_ _03074_ _03077_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07923__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09125__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13956_ _00287_ net101 clknet_leaf_56_clk DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_TAPCELL_ROW_17_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12907_ _02854_ _00397_ _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13887_ _00218_ net36 clknet_3_2__leaf_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_88_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12838_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-10\] _05723_ _05726_ _05727_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_97_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07439__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11235__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12769_ _05646_ _05650_ _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07197__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07611__A1 _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09980_ _02861_ _02862_ _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08931_ _06642_ _00382_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08862_ _00357_ _06674_ _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07813_ _00722_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08793_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-22\] _01608_ _01690_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07744_ net120 DDS_Stage.xPoints_Generator1.RegP\[-12\] _00684_ _00688_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09667__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07675_ _00641_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09414_ _02251_ _02303_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09345_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[11\] _02236_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_48_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_32_clk clknet_3_5__leaf_clk clknet_leaf_32_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_117_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09276_ _02084_ _02085_ _02166_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10985__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08227_ _01128_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07850__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08158_ _01058_ _01059_ _00954_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_30_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07109_ _06713_ _06645_ _06732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_120_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08089_ _00990_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08945__A4 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10120_ _02945_ _03001_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_98_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10051_ _02931_ _02933_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07905__A2 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09107__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13810_ _00141_ net36 clknet_leaf_52_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_145_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07343__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13741_ _00076_ net36 clknet_leaf_71_clk DDS_Stage.xPoints_Generator1.CosNew\[-12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_74_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10953_ _00381_ _00384_ _02499_ _02409_ _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_39_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13672_ _00007_ clknet_leaf_0_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10884_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[3\] _03674_ _03720_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[4\]
+ _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_128_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12623_ _03018_ _00378_ _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11217__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06892__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_23_clk clknet_3_6__leaf_clk clknet_leaf_23_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_155_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12554_ _04027_ _04028_ _05418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_136_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10976__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11505_ _04324_ _04346_ _04347_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10976__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07841__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12485_ _05339_ _05344_ _05345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11436_ _00378_ _01693_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11367_ _04209_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13106_ _05443_ _05832_ _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10318_ _03117_ _03120_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11940__A3 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11298_ _04121_ _04139_ _04140_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08149__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09346__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13037_ _05901_ _05939_ _05941_ _05942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10249_ _03044_ _03128_ _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11153__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09897__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10900__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11456__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13939_ _00270_ net101 clknet_leaf_31_clk net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07460_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-14\] _00472_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07391_ DDS_Stage.xPoints_Generator1.CosNew\[-2\] DDS_Stage.xPoints_Generator1.RegP\[-2\]
+ _00402_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_clk clknet_3_6__leaf_clk clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_29_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09130_ _02019_ _02022_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_151_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08085__A1 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08085__B2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ _01952_ _01954_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08012_ _06179_ _00388_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09034__B1 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08388__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09963_ _02838_ _02846_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08914_ _06664_ _00370_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09894_ _02697_ _02776_ _02777_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11144__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08845_ _01660_ _01661_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12892__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11695__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08560__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08776_ _01591_ _01671_ _01672_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07727_ _00678_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07658_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-7\] DDS_Stage.xPoints_Generator1.RegFrequency\[-7\]
+ _00626_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_67_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06874__A2 _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_7__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07589_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-4\] _05182_ _00570_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_36_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09328_ _02202_ _02218_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_146_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclone12 net141 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09812__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10958__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclone23 net146 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_63_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07823__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ _02150_ _02049_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclone56 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-19\] net155 vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlya_4
XFILLER_0_91_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12270_ _04953_ _04957_ _05113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11907__B1 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08379__A2 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11221_ _03817_ _03820_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_120_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11383__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07051__A2 _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11152_ _03340_ _00361_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10103_ _00388_ _06701_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_147_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11083_ _00372_ _02940_ _02938_ _00375_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10034_ _00373_ _06724_ _02807_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11985_ _04815_ _04827_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13724_ _00059_ net36 clknet_leaf_36_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_10936_ _03784_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10867_ _03706_ _03711_ _03737_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06865__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13655_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[0\] _06565_ _06608_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12606_ net84 _03558_ _05475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13586_ _03556_ _00397_ _06535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10798_ _03606_ _03607_ _03605_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_80_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12537_ _03018_ _00375_ _05400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12468_ _05017_ _05191_ _05209_ _05229_ _05327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_11419_ _00359_ _02236_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12399_ _04863_ _04864_ _05252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11374__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10177__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07042__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09319__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06960_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-19\] _06523_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xclkbuf_leaf_3_clk clknet_3_2__leaf_clk clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12874__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06891_ _05572_ _05442_ _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_08630_ _00428_ _01526_ _01527_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_55_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08561_ _06627_ _00379_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07512_ _05409_ _06458_ _00347_ _06753_ _05658_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08492_ _01390_ _01297_ _01391_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07443_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-17\] _00458_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13051__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07374_ _00407_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09113_ _06654_ _00382_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11601__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09044_ _01937_ _01913_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07281__A2 _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07033__A2 _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09946_ _00370_ _06730_ _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09877_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[17\] _02762_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09730__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09730__B2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08828_ _06649_ _00376_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_142_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_142_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _01581_ _01654_ _01655_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11770_ _04606_ _04611_ _04612_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_107_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10721_ _03584_ _03594_ _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_49_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13440_ _06300_ _06301_ _06376_ _06377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10652_ _03515_ _03518_ _03526_ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_76_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13371_ _06141_ _06285_ _06303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10583_ _03443_ _03458_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12322_ _05165_ _05166_ _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12253_ _05079_ _05094_ _05095_ _05096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13345__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10159__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_53_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11204_ _00390_ _02236_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07024__A2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12184_ _00397_ _01430_ _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XDDS_Module_41 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08772__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ _03972_ _03973_ _03976_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XDDS_Module_52 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_11066_ _03906_ _03907_ _03908_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA_clkbuf_leaf_68_clk_I clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09721__A1 _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10017_ _02896_ _02899_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11968_ _00359_ _02762_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07335__I0 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10095__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13707_ _00042_ clknet_leaf_39_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10919_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-12\] _03776_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11899_ _04741_ _04740_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_74_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10890__I0 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-25\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13638_ _06543_ _06548_ _06589_ _06590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10892__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13569_ _06454_ _06507_ _06515_ _06516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07090_ _05409_ _06715_ _06716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13336__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11347__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A2 _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09555__A4 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08763__A2 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09800_ _02593_ _02643_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07992_ _06642_ _00357_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07706__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09731_ _06664_ _00398_ _00394_ _06672_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06943_ _05420_ _05496_ _06340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09712__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09712__B2 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _02547_ _02548_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06874_ _05561_ _05583_ _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10322__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08613_ _01315_ _01322_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07869__A4 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09593_ _02480_ _02389_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_124_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08544_ _01373_ _01387_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12075__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08475_ _00379_ _06618_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10625__A3 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07426_ _05409_ _05984_ _06146_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07357_ _00396_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09876__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07288_ _05409_ _05702_ _05658_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_116_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09027_ _01840_ _01920_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_130_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11338__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07006__A2 _06623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10561__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09929_ _00388_ _00385_ _06691_ _06696_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_12940_ _05720_ _05722_ _05838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12871_ _05760_ _05666_ _05761_ _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07190__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11822_ _04660_ _04663_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13263__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07351__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11753_ _04594_ _04595_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_139_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10704_ net63 _06744_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11684_ _00372_ _01430_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08690__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10635_ _03037_ _03509_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13423_ _06358_ _06359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_153_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold68_I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13354_ _06223_ _06284_ _06285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10566_ _03432_ _03441_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07245__A2 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12305_ _05084_ _05085_ _05149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13318__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13285_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-5\] _06209_ _06210_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10497_ _03372_ _03373_ _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12236_ _00369_ _02236_ _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09537__A4 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10001__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10001__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12167_ _05007_ _05008_ _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_75_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11118_ _00397_ _02238_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12098_ _04938_ _04939_ _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11049_ _00372_ _02938_ _02854_ _00375_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput7 net133 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09170__A2 _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07181__A1 _06793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13730__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11265__B1 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11804__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08260_ _01155_ _01160_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07211_ _05409_ _06555_ _06787_ _06819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_117_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08191_ _01076_ _01092_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09225__A3 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07142_ _05409_ _05452_ _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_95_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09630__B1 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13797__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10240__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07073_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-2\] _06701_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11335__A4 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08200__A4 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07975_ _00842_ _00864_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09714_ _02520_ _02598_ _02599_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06926_ _06146_ _06114_ _06157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06857_ DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[3\] _05409_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_20
X_09645_ _02433_ _02434_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07172__A1 _06785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09576_ _02459_ _02463_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08527_ _01320_ _01426_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_104_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08458_ _01268_ _01269_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_34_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07475__A2 _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07409_ _06232_ _06645_ _05442_ _06146_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_80_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13548__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ _01287_ _01288_ _01289_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_107_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11559__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10420_ _03296_ _03297_ _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13788__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10351_ _03146_ _03228_ _03229_ _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06986__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13070_ _05952_ _05977_ _05978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_130_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10282_ _03160_ _03161_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12021_ _04164_ _04165_ _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13484__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07538__I0 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12923_ _05753_ _05818_ _05819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07163__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12039__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12854_ _05651_ _05718_ _05742_ _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06910__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11805_ _00361_ _01430_ _01249_ _00365_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12785_ _05663_ _05667_ _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_29_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09455__A3 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_1_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11736_ _04562_ _04578_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13539__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11667_ _04505_ _04506_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13406_ _06336_ _06339_ _06341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10618_ _03460_ _03465_ _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07218__A2 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11598_ _04425_ _04433_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11014__A3 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10549_ _03364_ _03367_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13337_ _06264_ _06266_ _06267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06977__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13268_ _06183_ _06192_ _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12219_ _05048_ _05060_ _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_90_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13199_ _06113_ _06117_ _06118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__10525__A2 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09391__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13951__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07760_ net4 DDS_Stage.xPoints_Generator1.RegP\[-4\] _00684_ _00696_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_108_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09143__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07691_ DDS_Stage.xPoints_Generator1.RegFrequency\[-3\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-3\]
+ _00650_ _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07154__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08497__A4 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09430_ _02310_ _02312_ _02318_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_121_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06901__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09361_ _02249_ _02250_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08312_ _01166_ _01168_ _01213_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09292_ _02092_ _02093_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_129_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08243_ _01137_ _01138_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08174_ _01043_ _01065_ _01075_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_119_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_119_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10213__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07125_ _06059_ _06668_ _06745_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08957__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06968__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07056_ _06059_ _06684_ _06686_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_132_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11308__A4 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13942__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13466__A1 _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07958_ _00858_ _00859_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09134__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06909_ _05442_ _05452_ _05973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07889_ net91 net142 net156 _06598_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07145__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09628_ _02426_ _02430_ _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09559_ _02378_ _02382_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12570_ _03971_ _04035_ _05436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_136_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09988__A4 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11521_ _04361_ _04362_ _04363_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_93_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11452_ net86 net83 _02409_ _02238_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_80_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10403_ _03037_ _03280_ _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_33_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11383_ net70 _01956_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06959__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10334_ _03204_ _03212_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13122_ net77 _06034_ _06035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_132_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13053_ _05878_ _05953_ _05959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_10265_ _03064_ _03143_ _03144_ _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11704__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12004_ _04786_ _04790_ _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_72_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08176__A3 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10196_ _02972_ _03075_ _03076_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13933__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08581__B1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07804__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09125__A2 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11468__B1 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13955_ _00286_ net101 clknet_leaf_56_clk DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_89_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12906_ _05798_ _05685_ _05799_ _05801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13886_ _00217_ net36 clknet_leaf_60_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_69_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12837_ _05623_ _05630_ _05725_ _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_69_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12768_ _05648_ _05649_ _05650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10443__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11719_ _00361_ _00365_ _01693_ _01610_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_51_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12699_ _05560_ _05575_ _05576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput10 net119 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08930_ _01730_ _01823_ _01824_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08861_ _01674_ _01755_ _01756_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13924__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07812_ _00376_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[23\] _00395_ _00722_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08792_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-22\] _01608_ _01689_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_74_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07714__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07743_ _00687_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07127__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07674_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-5\] _00640_ _00395_ _00641_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09413_ _02253_ _02302_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10682__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09344_ _05182_ _02234_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09275_ _00373_ _06674_ _02086_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_90_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08226_ net73 _05833_ _05398_ net60 _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10985__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09427__I0 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07850__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08157_ _00367_ _06308_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07108_ _06059_ _06729_ _06731_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ _06308_ _00355_ net152 net58 _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_3_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07039_ _05822_ _06672_ _06673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10050_ _02681_ _02932_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13915__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07624__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09107__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07118__A1 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12111__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_82_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13740_ _00075_ net36 clknet_leaf_69_clk DDS_Stage.xPoints_Generator1.CosNew\[-13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_138_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10952_ _00387_ _02238_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13671_ _00006_ clknet_leaf_77_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10883_ _03642_ _03733_ _03753_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_12622_ _05385_ _05490_ _05491_ _05492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10425__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12553_ _04027_ _04028_ _05417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_109_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10976__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11504_ _04326_ _04340_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_80_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07841__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12484_ _05343_ _05340_ _05344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_91_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12178__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11435_ _00372_ _01794_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11925__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11366_ _00390_ _01249_ _01247_ _00393_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_21_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ _03131_ _03152_ _03195_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13105_ _05830_ _05832_ _06016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11940__A4 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11297_ _04137_ _04138_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09346__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13036_ _05904_ _05920_ _05941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10248_ _03124_ _03127_ _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13906__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11153__A2 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10179_ _03056_ _03059_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10900__A2 _06777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07109__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12102__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08857__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13938_ _00269_ net101 clknet_leaf_31_clk net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_77_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13869_ _00200_ net36 clknet_leaf_54_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_76_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07390_ _00415_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07489__B _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08085__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09060_ _01796_ _01953_ _01873_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08011_ _06416_ _00382_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09034__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09034__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07596__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09962_ net55 _02839_ _02840_ _02845_ _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__10135__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08913_ _01805_ _01807_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_139_Left_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09893_ net61 net60 _06730_ _06738_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_110_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11144__A2 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08844_ _01664_ _01738_ _01739_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12892__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08775_ net61 net60 _06654_ _06659_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_97_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07726_ net110 DDS_Stage.xPoints_Generator1.RegF\[-5\] _00667_ _00678_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07657_ _00624_ _00625_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07520__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07588_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[27\] _00569_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10407__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09327_ _02204_ _02217_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_146_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone13 net141 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_118_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10958__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11080__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09258_ _02147_ _02148_ _02149_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone57 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-19\] net156 vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dlya_4
XFILLER_0_51_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08209_ _01099_ _01100_ _01110_ _01109_ _01108_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_09189_ _01918_ _02023_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11907__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11907__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11220_ _04058_ _04061_ _04062_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08379__A3 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07587__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11383__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11151_ _00369_ _03189_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10102_ _00382_ _06710_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11082_ _00372_ _00375_ _02940_ _02938_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_147_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10033_ _02801_ _02914_ _02915_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10894__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11984_ _04819_ _04826_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13723_ _00058_ net36 clknet_leaf_21_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10935_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-4\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-4\]
+ _05171_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_27_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07511__A1 _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13654_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[0\] _06565_ _06567_ _06607_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10866_ _03704_ _03712_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12605_ _03556_ _00359_ _05473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13585_ _06482_ _06474_ _06533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10797_ _03668_ _03669_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12536_ _02940_ _00378_ _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_81_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12467_ _05319_ _05323_ _05325_ _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_152_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11418_ net87 _02409_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12398_ _04869_ _05251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11374__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11349_ _04190_ _04191_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09319__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13019_ _05863_ _05922_ _05923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06890_ _05409_ _05529_ _05658_ _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12874__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08560_ _06637_ _00373_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07511_ _06703_ _06629_ _06766_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08491_ _01278_ _01291_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11834__B1 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07442_ _05409_ _05973_ _06622_ _06816_ _00456_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07373_ DDS_Stage.xPoints_Generator1.CosNew\[-11\] DDS_Stage.xPoints_Generator1.RegP\[-11\]
+ _00402_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08058__A2 _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13051__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09112_ _01905_ _02003_ _02004_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09043_ _01921_ _01923_ _01936_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_147_Left_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09945_ _02826_ _02828_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_5_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09876_ _02681_ _02759_ _05182_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09730__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08827_ _06642_ _00379_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_142_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ _01583_ _01596_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10628__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_156_Left_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07709_ _00669_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08689_ _01584_ _01585_ _01586_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_138_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10720_ _03586_ _03593_ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_24_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10651_ _03311_ _03525_ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10582_ _03446_ _03449_ _03457_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13370_ _06300_ _06301_ _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12321_ _05158_ _05159_ _05166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12252_ _05080_ _05081_ _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_133_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11203_ _00397_ _02051_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12183_ _05020_ _05025_ _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11134_ _03972_ _03973_ _03976_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XDDS_Module_42 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_11065_ net54 _03340_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10016_ _02897_ _02898_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09721__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07812__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11967_ _00354_ _02854_ _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07335__I1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13706_ _00041_ clknet_3_5__leaf_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10095__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10918_ _03775_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11898_ _04464_ _04465_ _04413_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_156_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13637_ _06539_ _06549_ _06589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10849_ _00552_ _03720_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13568_ _06457_ _06506_ _06515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12519_ _03485_ _00359_ _05380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07263__A3 _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13499_ _06438_ _06440_ _06441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11347__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07991_ _00852_ _00891_ _00892_ _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09730_ _06664_ _00398_ _00394_ _06672_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06942_ _06059_ _06297_ _06319_ _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10858__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09712__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09661_ _00376_ _06696_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06873_ _05572_ _05474_ _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_119_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08612_ _01314_ _01323_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_94_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09592_ _02327_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_124_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07722__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08543_ _01363_ _01419_ _01441_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08474_ _06633_ _00373_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07425_ _05420_ _06092_ _05561_ _06232_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__09228__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07356_ _00393_ _00394_ _00395_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12783__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07287_ _00295_ _00341_ _06146_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_131_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09026_ _01916_ _01919_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11338__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10561__A3 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ _00382_ _06701_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10849__A1 _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09859_ _02741_ _02743_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12870_ net66 net54 _03725_ _03727_ _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07190__A2 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07632__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11821_ _04660_ _04663_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13263__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11274__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11752_ _04498_ _04499_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_64_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10703_ _03115_ _03576_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11683_ _00378_ _01247_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__A2 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11026__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13422_ _06316_ _06357_ _06358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10634_ net57 _02704_ _03508_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07587__B _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13353_ _06231_ _06283_ _06284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10565_ _03373_ _03440_ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12304_ _04371_ _04385_ _05147_ _05148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13284_ _06204_ _06208_ _06209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10496_ _00398_ _00394_ _06710_ _06724_ _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_121_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12526__A1 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12235_ _05077_ _05074_ _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10001__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12166_ _05007_ _05008_ _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_75_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11117_ _03955_ _03959_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12097_ _04938_ _04939_ _04940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11048_ _00372_ _00375_ _02938_ _02854_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xinput8 net131 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09458__A1 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12999_ _05806_ _05815_ _05900_ _05901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11265__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11265__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07210_ _06818_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11017__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08190_ _01083_ _01091_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07141_ _05431_ _06759_ _05420_ _06760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09225__A4 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09630__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09630__B2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07072_ _05658_ _06699_ _06700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12517__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08197__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ _00874_ _00875_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09713_ net91 net143 _06710_ _06724_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06925_ _05647_ _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_20
X_09644_ _02433_ _02434_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06856_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-25\] _05398_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_93_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09575_ _02460_ _02461_ _02462_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_78_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08526_ _00424_ _01349_ _01425_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_148_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_52_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08457_ _01258_ _01355_ _01356_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07408_ _05409_ _05474_ _05518_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08388_ net96 _06179_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11559__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_67_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07339_ _00381_ _00382_ _05182_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10350_ _03147_ _03148_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_60_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06986__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09009_ _01827_ _01828_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10281_ _03155_ _03156_ _03159_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_103_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13181__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12020_ net89 _04857_ _04862_ _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__13484__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12922_ _05794_ _05817_ _05818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07163__A2 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12853_ _05654_ _05717_ _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11804_ _00369_ _01247_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12784_ _05664_ _05665_ _05666_ _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_29_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09455__A4 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11735_ _04561_ _04562_ _04563_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09860__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11666_ _04508_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13405_ _06337_ _06338_ _06339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10617_ _03424_ _03459_ _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08415__A2 _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09612__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11597_ _04420_ _04438_ _04439_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__11014__A4 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13336_ net147 _00390_ _06266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10548_ _03378_ _03394_ _03423_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13267_ _06186_ _06191_ _06192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10479_ _03274_ _03314_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08179__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13172__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12218_ _05048_ _05060_ _05061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_90_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13198_ _06014_ _06115_ _06116_ _06117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07926__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12149_ net66 net54 _02586_ net135 _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07690_ DDS_Stage.xPoints_Generator1.RegFrequency\[-3\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-3\]
+ _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06901__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _00370_ _06691_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08103__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08311_ _01170_ _01194_ _01197_ _01212_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XPHY_EDGE_ROW_111_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09291_ _02178_ _02181_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08242_ _01121_ _01142_ _01143_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_145_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08173_ _01047_ _01064_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_119_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_119_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07124_ _05280_ _06744_ _06745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06968__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07090__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07055_ _05822_ _06685_ _06686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09906__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_120_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07957_ _06649_ net138 _00391_ _05833_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06908_ _05409_ _05442_ _05875_ _05930_ _05951_ _05962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_07888_ net91 net156 _06598_ net142 _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_39_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07145__A2 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-24\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09627_ _02437_ _02445_ _02513_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06839_ _05182_ net18 _05193_ _05204_ _05215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_78_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09558_ _02421_ _02437_ _02445_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__12977__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08509_ _01282_ _01407_ _01408_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09489_ _02267_ _02376_ _02377_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11520_ _00359_ _02409_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12729__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11451_ net86 _02409_ _02238_ net83 _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10402_ _02608_ _02704_ _03279_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_132_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11382_ _04175_ _04223_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_59_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06959__A2 _06502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13121_ _05842_ _05933_ _06034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10333_ _03126_ _03211_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13052_ _05955_ _05956_ _05957_ _05958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_103_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10264_ _03065_ _03066_ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11704__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12003_ _04802_ _04844_ _04845_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_72_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08176__A4 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10195_ _02975_ _02989_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_100_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08581__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08581__B2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11468__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13954_ _00285_ net36 clknet_leaf_59_clk DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09125__A3 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11468__B2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07136__A2 _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12905_ _05687_ _05799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_17_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13885_ _00216_ net36 clknet_leaf_55_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_115_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12836_ _05619_ _05622_ _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_97_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12767_ _02586_ _00397_ _05601_ _05649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08636__A2 _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11718_ _00369_ _01524_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12698_ _05569_ _05574_ _05575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 net117 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11649_ _04488_ _04491_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_154_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13319_ _06245_ _06246_ _06247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07072__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13145__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08860_ net61 net60 _06664_ _06659_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_07811_ _00721_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08791_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-21\] _01614_ _01687_ _01688_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_74_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07742_ net114 DDS_Stage.xPoints_Generator1.RegP\[-13\] _00684_ _00687_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11459__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07673_ DDS_Stage.xPoints_Generator1.CosNew\[-5\] _00639_ _00577_ _00640_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09412_ _02273_ _02301_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10682__A2 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08088__B1 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09343_ _02229_ _02232_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_101_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09824__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10434__A2 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11631__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09274_ _02079_ _02097_ _02164_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08225_ _01125_ _01126_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_90_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13860__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09427__I1 _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08156_ _00363_ _06416_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11395__B1 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07063__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07107_ _05822_ _06730_ _06731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08087_ net58 _06308_ _00355_ net152 _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_101_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07038_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-8\] _06672_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_2_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11698__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08989_ _01817_ _01831_ _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_145_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07118__A2 _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12111__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10951_ _00397_ _02236_ _03793_ _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_138_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06877__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13670_ _00005_ clknet_leaf_78_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10882_ _03736_ _03738_ _03752_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_78_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12621_ _05386_ _05388_ _05491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_38_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10425__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12552_ _05412_ _05415_ _05416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11503_ _04326_ _04340_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_109_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13851__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12483_ _05342_ _05343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_22_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12178__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11434_ _00375_ _01792_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11925__A2 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11365_ _04194_ _04206_ _04207_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13104_ _06014_ _06015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_120_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10316_ _03114_ _03130_ _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11296_ _04137_ _04138_ _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13035_ _05904_ _05920_ _05939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10247_ _03125_ _03126_ _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11689__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10178_ _03057_ _03058_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07109__A2 _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12102__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13937_ _00268_ net101 clknet_3_5__leaf_clk net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_44_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08857__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06868__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13868_ _00199_ net36 clknet_leaf_65_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12819_ _05608_ _05609_ _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_146_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13799_ _00130_ net36 clknet_leaf_60_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[27\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_84_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07489__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07293__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08010_ _00832_ _00911_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_71_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13366__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09034__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07045__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09961_ _02842_ _02843_ _02844_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_111_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08912_ _01723_ _01724_ _01806_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09892_ net61 _06730_ _06738_ net60 _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11144__A3 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08843_ _01666_ _01679_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10352__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08774_ net61 _06654_ _06659_ net60 _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07725_ _00677_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10104__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07656_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-8\] DDS_Stage.xPoints_Generator1.RegFrequency\[-8\]
+ _00620_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07587_ _05387_ _00567_ _00568_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09326_ _02212_ _02216_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11604__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07399__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclone14 net67 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XANTENNA__07284__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09257_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-17\] _02149_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11080__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone36 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[15\] net135 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_4
XFILLER_0_90_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08208_ _01108_ _01109_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09188_ _02019_ _02022_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11907__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07036__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08139_ _05398_ _00379_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08379__A4 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13109__A1 _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11150_ _03988_ _03992_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10101_ _02903_ _02981_ _02982_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_8_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11081_ _03923_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_147_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08536__B2 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10032_ _02803_ _02819_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10343__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10894__A2 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-23\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11983_ _04822_ _04825_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13722_ _00057_ clknet_leaf_15_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11843__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10934_ _03783_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07511__A2 _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13653_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[1\] _06573_ _06605_ _06606_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10865_ _03688_ _03734_ _03735_ _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_151_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13596__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12604_ _05380_ _05470_ _05471_ _05472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13584_ _06488_ _06497_ _06531_ _06532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10796_ _03560_ _03604_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_80_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07275__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12535_ _03994_ _05395_ _05396_ _05397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12466_ _03768_ _05321_ _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07027__A1 _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11417_ net84 _02238_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08224__B1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12397_ _04742_ _05230_ _05241_ _05249_ _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_151_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08775__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11348_ _00372_ _01693_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11279_ _00372_ _00375_ _02584_ _02499_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_13018_ _05898_ _05921_ _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12874__A3 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07510_ _00510_ _00511_ _00512_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08490_ _01278_ _01291_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11834__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11834__B2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07441_ _06146_ _05463_ _06125_ _00455_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_119_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13587__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07372_ _00406_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09111_ _01906_ _01907_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13815__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07266__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _01927_ _01935_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_98_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07018__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09944_ _02723_ _02724_ _02827_ _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_5_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09875_ _02681_ _02759_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09191__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08826_ _06654_ _00373_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12078__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08757_ _01583_ _01596_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07708_ net8 DDS_Stage.xPoints_Generator1.RegF\[-14\] _00667_ _00669_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10628__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08688_ net95 net155 _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_107_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07639_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-10\] _00610_ _00395_ _00611_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10650_ _03521_ _03524_ _03525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_137_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13806__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07257__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09309_ _06642_ _06637_ _00398_ _00394_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_36_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10581_ _03311_ _03456_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_62_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12320_ _05140_ _05144_ _05165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07009__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12251_ _05080_ _05081_ _05094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10939__I0 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11202_ _04043_ _04044_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07804__I0 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12182_ _05021_ _05024_ _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11133_ _03950_ _03974_ _03975_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XDDS_Module_43 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__07365__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11064_ net87 _03416_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09182__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10015_ _00376_ _06724_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11816__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11966_ _00351_ _02938_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_82_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13705_ _00040_ clknet_leaf_34_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10917_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-13\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-13\]
+ _05171_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07496__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11897_ _04413_ _04516_ _04736_ _04739_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_74_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13636_ _00390_ _03725_ _06588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10848_ _03683_ _03719_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07248__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13567_ _05822_ _06512_ _06514_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10779_ _03636_ _03651_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12518_ _03989_ _05377_ _05378_ _05379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13498_ _06439_ _06372_ _06440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12449_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-24\] _05300_ _05306_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10555__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_93_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07420__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07990_ net91 _00363_ _06633_ _06627_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_120_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06941_ _05822_ _06308_ _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09660_ _00379_ _06691_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06872_ _05420_ _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_16
XFILLER_0_94_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08611_ _01509_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09591_ _02414_ _02478_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_124_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08542_ _01366_ _01418_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_124_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07487__A1 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08473_ _00885_ _01296_ _01372_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07424_ _06630_ _00441_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09228__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07239__A1 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07355_ _05171_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XANTENNA__12232__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone10_I net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12783__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07286_ _05583_ _06711_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09025_ _01917_ _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07411__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10561__A4 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09927_ _02730_ _02809_ _02810_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09858_ _02629_ _02630_ _02742_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08911__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08809_ _01632_ _01682_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09789_ _02048_ _02145_ _02397_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_11820_ _04661_ _04662_ _04625_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_96_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11751_ _04574_ _04582_ _04593_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_64_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07478__A1 _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11274__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _03037_ _03509_ _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11682_ _04521_ _04524_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_126_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13421_ _06318_ _06356_ _06357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_138_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10633_ net63 _06742_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11026__A2 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13352_ _06234_ _06282_ _06283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10564_ _03435_ _03439_ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_134_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12303_ _04357_ _04370_ _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_51_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13283_ _06015_ _06026_ _06113_ _06207_ _06208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_10495_ _00398_ _06710_ _06724_ _00394_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12234_ _05075_ _05076_ _04990_ _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__12526__A2 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12165_ _04914_ _04932_ _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11116_ _03956_ _03957_ _03958_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_12096_ _04801_ _04859_ _04939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11047_ _03889_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput9 net113 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_24_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09458__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12998_ _05809_ _05899_ _05900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07469__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11265__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11949_ _04779_ _04791_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_71_clk clknet_3_0__leaf_clk clknet_leaf_71_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12214__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11017__A2 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13619_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[0\] _06565_ _06569_ _06570_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_55_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07140_ _06232_ _05463_ _06759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09630__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07071_ _05409_ _05485_ _05507_ _06698_ _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_33_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12517__A2 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08197__A2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07973_ _06627_ _00370_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09712_ net91 _06710_ _06724_ net143 _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06924_ _05658_ _06125_ _06135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09643_ _02516_ _02529_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06855_ _05171_ _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ _00385_ _06674_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08525_ _01422_ _01424_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_78_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_62_clk clknet_3_3__leaf_clk clknet_leaf_62_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_46_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _01259_ _01272_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_46_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07407_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-23\] _00428_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08387_ _00352_ _06659_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07338_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-6\] _00382_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
XFILLER_0_61_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07269_ _05409_ _05485_ _05561_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_131_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ _01827_ _01828_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_150_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10280_ _03155_ _03156_ _03159_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13181__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12921_ _05797_ _05801_ _05816_ _05817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_88_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12852_ _05648_ _05649_ _05646_ _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_38_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11803_ _00361_ _00365_ _01430_ _01249_ _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_12783_ net70 _03679_ _05666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_53_clk clknet_3_1__leaf_clk clknet_leaf_53_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11734_ _04575_ _04529_ _04576_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_84_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09860__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11665_ _04482_ _04483_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10616_ _03401_ _03463_ _03490_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13404_ _03485_ _00390_ _06338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ _04435_ _04437_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09612__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13335_ _03340_ _00393_ _06264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10547_ _03362_ _03377_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13266_ _06187_ _06188_ _06189_ _06191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10478_ _03353_ _03354_ _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08179__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13172__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12217_ _05055_ _05059_ _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_90_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13197_ _06008_ _06013_ _06116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_90_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11183__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07926__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12148_ net66 _02586_ net135 net54 _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09128__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12079_ _00354_ _02762_ _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_44_clk clknet_3_4__leaf_clk clknet_leaf_44_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08103__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _01177_ _01199_ _01211_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_59_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09290_ _02179_ _02180_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10997__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08241_ _01119_ _01120_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_31_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08172_ _01072_ _01073_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07123_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[5\] _06744_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_119_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07728__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07054_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-5\] _06685_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_88_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_132_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07956_ _06649_ _00352_ _00391_ _05833_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06907_ _05474_ _05940_ _05951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07887_ _00787_ _00788_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06838_ DDS_Stage.LCU.state\[2\] DDS_Stage.LCU.state\[0\] DDS_Stage.LCU.state\[1\]
+ _05204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09626_ _02423_ _02436_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09557_ _02438_ _02441_ _02444_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_78_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ _06642_ net61 net60 _06637_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__12977__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09488_ _02268_ _02269_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_148_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10988__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08439_ _01221_ _01222_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_93_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11450_ _04264_ _04268_ _04292_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12729__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10401_ net63 _06724_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11381_ _04175_ _04223_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_34_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07638__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13120_ _05847_ _06031_ _06032_ _06033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_150_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10332_ _03207_ _03210_ _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13051_ _00361_ _03727_ _05957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10263_ _03065_ _03066_ _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_108_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12002_ _04830_ _04843_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_72_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10194_ _02975_ _02989_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10912__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08581__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07373__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11468__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13953_ _00284_ net36 clknet_leaf_58_clk DDS_Stage.Block_Cosine.PolyRAM_1.MEM_A0.addr\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__09125__A4 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12904_ _05681_ _05798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13884_ _00215_ net36 clknet_leaf_59_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_17_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12835_ _05720_ _05722_ _05723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclkbuf_leaf_26_clk clknet_3_7__leaf_clk clknet_leaf_26_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08097__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12766_ _05599_ _05600_ _05648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_127_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10979__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11717_ _04556_ _04559_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12697_ _05570_ _05571_ _05573_ _05574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_25_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11648_ _04489_ _04490_ _04443_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
Xinput12 net111 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11579_ _00372_ _00375_ _01610_ _01524_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_25_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13318_ _00372_ _03727_ _06246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13145__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13249_ _06099_ _06172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07810_ _00373_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[22\] _00395_ _00721_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08790_ _01616_ _01686_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07741_ _00686_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11459__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_66_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09521__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07672_ DDS_Stage.xPoints_Generator1.RegFrequency\[-5\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-5\]
+ _00638_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_36_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09411_ _02275_ _02300_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_clk clknet_3_7__leaf_clk clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09342_ _02229_ _02232_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08088__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08088__B2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09824__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09273_ _02082_ _02096_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_8_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11631__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08224_ net58 _06179_ _05864_ _00355_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_106_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11919__B1 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08155_ _01031_ _01055_ _01056_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11395__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11395__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07106_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[2\] _06730_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_28_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08086_ _00987_ _00982_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_140_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07037_ _06667_ _06670_ _06671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_19_clk_I clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11147__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08012__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11698__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08988_ _01817_ _01831_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07193__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07939_ _00803_ _00817_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12647__A1 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10950_ _03790_ _03791_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09609_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-13\] _02394_ _02406_ _02497_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10881_ _03082_ _03741_ _03751_ _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06877__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12620_ _05386_ _05388_ _05490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07826__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12551_ _05413_ _05414_ _05415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11083__B1 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11502_ _04225_ _04343_ _04344_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_53_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12482_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-17\] _05341_ _05342_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11433_ _04246_ _04274_ _04275_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11364_ _04200_ _04205_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10315_ _03192_ _03193_ _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13103_ _06008_ _06013_ _06014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11295_ _04045_ _04049_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13034_ _05861_ _05923_ _05937_ _05938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10246_ _00398_ _00394_ _06696_ _06701_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_120_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11689__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09751__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10177_ _00376_ _06738_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12638__A1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13936_ _00267_ net101 clknet_leaf_16_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11310__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06868__A2 _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13867_ _00198_ net36 clknet_3_0__leaf_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_TAPCELL_ROW_85_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13063__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12818_ _05700_ _05704_ _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13798_ _00129_ net36 clknet_leaf_64_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[26\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_139_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12749_ _05623_ _05630_ _05631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_41_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_116_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09990__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09960_ _02841_ _02753_ _02756_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_6_clk clknet_3_3__leaf_clk clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08911_ _06654_ _00373_ _01725_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09891_ _02701_ _02705_ _02774_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09742__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08842_ _01666_ _01679_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11144__A4 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10352__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08773_ _01667_ _01668_ _01669_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07724_ net106 DDS_Stage.xPoints_Generator1.RegF\[-6\] _00667_ _00677_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07356__I0 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10104__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07655_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-8\] DDS_Stage.xPoints_Generator1.RegFrequency\[-8\]
+ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07586_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-5\] _05182_ _00568_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09325_ _02213_ _02214_ _02215_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_75_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11604__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09256_ _01969_ _01973_ _02047_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone48 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[25\] net147 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_4
X_08207_ _00992_ _01001_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_7_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclone59 net159 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09187_ _02002_ _02010_ _02078_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07188__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08138_ _05833_ _00376_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08069_ _00948_ _00969_ _00970_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10100_ _02904_ _02905_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11080_ _00378_ _02854_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10031_ _02803_ _02819_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10343__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11982_ _04823_ _04824_ _04149_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__07347__I0 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13721_ _00056_ clknet_leaf_20_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10933_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-5\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-5\]
+ _05171_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11843__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10864_ _03690_ _03715_ _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13652_ _06575_ _06579_ _06604_ _06605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_128_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12603_ _03556_ net66 net54 _03558_ _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_66_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13596__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10795_ _03563_ _03603_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13583_ _06492_ _06530_ _06531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07275__A2 _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12534_ _03995_ _03996_ _05396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_35_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12465_ _03768_ _05321_ _05322_ _05323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_124_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11359__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08224__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11416_ _04243_ _04257_ _04258_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07027__A2 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12396_ _05244_ _05247_ _05229_ _05017_ _05249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__08224__B2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11347_ _00375_ _01610_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08775__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09972__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12859__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11278_ _04111_ _04114_ _04120_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13017_ _05901_ _05904_ _05920_ _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10229_ _03072_ _03083_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13919_ _00250_ net36 clknet_leaf_34_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11834__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07440_ _06232_ _05940_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_58_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13587__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07371_ DDS_Stage.xPoints_Generator1.CosNew\[-12\] DDS_Stage.xPoints_Generator1.RegP\[-12\]
+ _00402_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09110_ _01906_ _01907_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_128_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09041_ _01930_ _01934_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_26_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07018__A2 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10022__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09943_ _00373_ _06710_ _02725_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09715__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09874_ _02758_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09191__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08825_ _01719_ _01720_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13751__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12078__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ _01634_ _01652_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_142_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07707_ _00668_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10628__A3 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08687_ net137 _06674_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07638_ DDS_Stage.xPoints_Generator1.CosNew\[-10\] _00609_ _00577_ _00610_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_24_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07569_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[18\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\]
+ _00395_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09308_ _06637_ _00398_ _00394_ _06642_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_152_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10580_ _03452_ _03455_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _02130_ _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12250_ _05042_ _05092_ _05093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12002__A2 _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11201_ _03795_ _03798_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10013__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12181_ _05022_ _05023_ _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07646__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11132_ _03952_ _03966_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_101_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_79_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XDDS_Module_44 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_101_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11063_ _00359_ _03266_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10014_ _00379_ _06710_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09182__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13742__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07381__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11965_ _04805_ _04806_ _04807_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11816__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_82_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13704_ _00039_ clknet_leaf_39_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10916_ _05387_ _03773_ _03774_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08693__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07496__A2 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11896_ _04737_ _04738_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_88_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13635_ _00393_ _03679_ _06586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10847_ _03717_ _03718_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13566_ _05280_ net24 _06514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10778_ _03639_ _03650_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12517_ _03556_ net86 net83 _03485_ _05378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_13497_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-3\] _06364_ _06439_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12448_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-24\] _05300_ _05304_ _05305_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12379_ _05017_ _05191_ _05209_ _05229_ _05230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_1_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_97_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06940_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-21\] _06308_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07355__I _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06871_ _05420_ _05550_ _05561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13733__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08610_ _01422_ _01424_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09590_ _02416_ _02477_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13257__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06931__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08541_ _01438_ _01439_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_124_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08472_ _01293_ _01370_ _01371_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_106_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07423_ _05778_ _06754_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-2\] _00394_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_0_9_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12232__A2 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10243__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07285_ _00339_ _00340_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06998__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09024_ _00398_ _00394_ _06627_ _06618_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07798__I0 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07947__B1 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09926_ _02731_ _02732_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13496__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09857_ _00373_ _06708_ _02631_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07175__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13724__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08808_ _01702_ _01703_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08911__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06922__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09788_ _02399_ _02403_ _02672_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06922__B2 _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08739_ _01481_ _01580_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08124__B1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11750_ _04572_ _04573_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_64_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10701_ _03503_ _03574_ _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_37_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11681_ _04522_ _04521_ _04523_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_83_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13420_ _06331_ _06355_ _06356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10632_ _03115_ _03506_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10563_ _03436_ _03438_ _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13351_ _06256_ _06281_ _06282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06989__A1 _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12302_ _05145_ _05146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10494_ _02704_ _03369_ _03370_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13282_ _06116_ _06205_ _06206_ _06207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12233_ _00351_ _02586_ _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12164_ _04987_ _05005_ _05006_ _05007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_3_0__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11115_ _02762_ _00381_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12095_ _04913_ _04936_ _04937_ _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11046_ _00378_ _02762_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07166__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06913__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12997_ _05814_ _05899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_86_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11948_ _04786_ _04790_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08666__A1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07469__A2 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11879_ _04686_ _04720_ _04721_ _04714_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_74_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13618_ _06568_ _06511_ _06569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12214__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13549_ _00387_ _03679_ _06495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11973__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07070_ _05409_ _06340_ _06698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_70_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12517__A3 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13954__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07972_ _00870_ _00873_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09711_ _02524_ _02528_ _02596_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06923_ _05572_ _05442_ _06125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__07157__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09642_ _02524_ _02528_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06854_ _05366_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06904__A1 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09573_ _00388_ _06672_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08524_ _01251_ _01309_ _01423_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_148_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10464__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08455_ _01273_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_46_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07406_ _05387_ _00424_ _00427_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08386_ _06654_ _00355_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13402__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07337_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-6\] _00381_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_0_151_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__A2 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11964__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07268_ _06232_ _06125_ _06727_ _06753_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_143_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09007_ _01897_ _01900_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_150_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07199_ _05182_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-16\] _06810_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07396__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13945__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09909_ _02791_ _02792_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12920_ _05806_ _05815_ _05816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12851_ _05636_ _05733_ _05735_ _05360_ _05739_ _05740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_68_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11802_ _04623_ _04639_ _04640_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_68_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12782_ net86 _03727_ _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11733_ _04527_ _04528_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11664_ _04505_ _04506_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13403_ net147 _00393_ _06337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10615_ _03082_ _03464_ _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11595_ _04435_ _04437_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_153_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13334_ _03266_ _00397_ _06263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10546_ _03420_ _03421_ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13265_ _03556_ _00381_ _06189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10477_ _03082_ _03320_ _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12216_ _05056_ _05057_ _05058_ _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_20_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13196_ _05829_ _05840_ _05928_ _06024_ _05927_ _06115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_121_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13936__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_90_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11183__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07926__A3 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12147_ _00359_ _02499_ _04990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09128__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12078_ _00351_ _02854_ _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13782__D _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11029_ net66 net54 _03266_ _03189_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10694__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08103__A3 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11643__B1 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08240_ _01140_ _01141_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10997__A2 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12199__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08171_ _06308_ _00370_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_83_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09064__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11946__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07122_ _06059_ _06741_ _06743_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_119_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _06146_ _06683_ _06684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13927__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07744__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07955_ _06642_ _00355_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12123__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06906_ _05420_ _05431_ _05940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07886_ _06637_ net58 _00355_ _06633_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_39_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10685__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09625_ _02421_ _02510_ _02511_ _02446_ _02467_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_06837_ net17 _05193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07550__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09556_ _02442_ _02443_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08507_ _06642_ net60 _06637_ net61 _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09487_ _02268_ _02269_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10988__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08438_ _00945_ _00978_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_92_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08369_ _01268_ _01269_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11937__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10400_ _03115_ _03277_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11380_ _04187_ _04221_ _04222_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_22_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10331_ _03208_ _03209_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_132_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13050_ _00365_ _03725_ _05956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10262_ _03138_ _03141_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13918__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12001_ _04830_ _04843_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_44_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10193_ _00373_ _06738_ _02979_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13952_ _00283_ net101 clknet_leaf_26_clk net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_12903_ _05705_ _05714_ _05796_ _05797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13883_ _00214_ net36 clknet_leaf_60_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07541__A1 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12834_ _05544_ _05618_ _05721_ _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_87_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08097__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12765_ _05595_ _05644_ _05645_ _05646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_68_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10979__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11716_ _04557_ _04558_ _04485_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_126_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12696_ _03556_ _00361_ _05573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11647_ net66 _02051_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput13 net115 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11578_ _00378_ _01430_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13317_ _00375_ _03725_ _06245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10600__A1 _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10529_ _03272_ _03322_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13248_ _06149_ _06170_ _06171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_0_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13909__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13179_ _03340_ _00387_ _06096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07740_ net8 DDS_Stage.xPoints_Generator1.RegP\[-14\] _00684_ _00686_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09521__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ _00636_ _00637_ _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09410_ _02291_ _02299_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09809__B1 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ _02150_ _02049_ _02230_ _02231_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_87_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08088__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09824__A3 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11092__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09272_ _02075_ _02129_ _02162_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_47_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08223_ net58 _00355_ _06179_ _05864_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_56_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09037__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11919__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11919__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08154_ net91 net142 _06308_ _06179_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_67_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07599__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11395__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12592__A1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07105_ _06146_ _06728_ _06729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08085_ _05398_ _00376_ _00373_ _05833_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_141_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07036_ _05658_ _05680_ _06669_ _06670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11147__A2 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08012__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08987_ _01810_ _01879_ _01880_ _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_138_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07938_ _00837_ _00839_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__12647__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10658__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07869_ net137 _00355_ _06633_ _06627_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_3_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09608_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-12\] _02495_ _02496_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_10880_ _03743_ _03745_ _03750_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09539_ _00357_ _06724_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_51_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11083__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12550_ _02586_ _00390_ _05414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07826__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11083__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11501_ _04289_ _04342_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12481_ _05336_ _05268_ _05341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11432_ _04247_ _04248_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_22_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12583__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11363_ _04200_ _04205_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13102_ _06010_ _06012_ _06013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10314_ _03154_ _03163_ _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_60_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_131_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11294_ _04127_ _04135_ _04136_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13033_ _05863_ _05922_ _05937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10245_ _00398_ _06696_ _06701_ _00394_ _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09200__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10897__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10176_ _00379_ _06730_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09751__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12638__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10649__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13935_ _00266_ net101 clknet_leaf_20_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11310__A2 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13866_ _00197_ net36 clknet_leaf_74_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_TAPCELL_ROW_85_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12817_ _05701_ _05703_ _05704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13063__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13797_ _00128_ net36 clknet_leaf_50_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_57_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12748_ _05445_ _05626_ _05629_ _05630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_45_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12679_ _05549_ _05553_ _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_41_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09990__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12326__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08910_ _01718_ _01736_ _01804_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09890_ _02696_ _02700_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07202__B1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08841_ _01718_ _01736_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09742__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08772_ net95 _06598_ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07723_ _00676_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_108_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07505__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07356__I1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07654_ _00623_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07585_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[26\] _00567_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11065__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09324_ _06649_ net95 _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09255_ _01968_ _01961_ _02146_ _02057_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_146_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone38 net140 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_91_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08206_ _01101_ _01106_ _01107_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_44_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09186_ _02005_ _02009_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08137_ _05864_ _00373_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08068_ _00967_ _00968_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13711__CLK clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07992__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07019_ _06059_ _06653_ _06655_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_147_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10030_ _02864_ _02912_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_126_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11981_ _00354_ _02938_ _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07347__I1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13720_ _00055_ clknet_leaf_16_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10932_ _05822_ _00312_ _03782_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_27_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13651_ _06581_ _06584_ _06603_ _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_67_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10863_ _03690_ _03715_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12602_ _03556_ net54 _03558_ net66 _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11056__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13582_ _06496_ _06530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_50_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10794_ _03629_ _03632_ _03666_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_67_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12533_ _03995_ _03996_ _05395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_135_Left_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_80_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07379__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12464_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-19\] _05317_ _05322_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11359__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12556__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_65_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11415_ net66 net54 _02238_ _02236_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_62_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12395_ _05245_ _05246_ _05247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08224__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11346_ _04188_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08775__A3 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11277_ _04115_ _04119_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12859__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13016_ _05910_ _05918_ _05920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09724__A2 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _03027_ _03071_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10159_ net63 _06696_ _02608_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13284__A2 _06208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13918_ _00249_ net36 clknet_leaf_39_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-17\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_89_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13849_ _00180_ net36 clknet_leaf_69_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_57_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_18_clk_I clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07370_ _00405_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09660__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09040_ _01931_ _01932_ _01933_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_154_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10022__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09942_ _02825_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09715__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09873_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-9\] _02755_ _02757_ _02758_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_110_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ _01578_ _01663_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07752__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08755_ _01637_ _01651_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_142_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07706_ net2 DDS_Stage.xPoints_Generator1.RegF\[-15\] _00667_ _00668_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11286__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08686_ _00355_ _06672_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10628__A4 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07637_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-10\] DDS_Stage.xPoints_Generator1.RegFrequency\[-10\]
+ _00608_ _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_24_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07568_ _00558_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12786__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09307_ _02112_ _02196_ _02197_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_118_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07499_ _05171_ _00503_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09238_ _02075_ _02129_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12538__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09169_ _01695_ _01698_ _02053_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09403__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11200_ _04042_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11210__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10013__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12180_ _00381_ _01794_ _01792_ _00384_ _05023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09954__A2 _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11131_ _03952_ _03966_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDDS_Module_45 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_11062_ _03874_ _03903_ _03904_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10013_ _00373_ _06730_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11964_ net66 net83 _02854_ _02762_ _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_98_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11816__A3 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08142__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13703_ _00038_ clknet_leaf_47_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10915_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-14\] _03774_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11895_ _04513_ _04514_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08693__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07496__A3 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11029__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13634_ _06557_ _06558_ _06556_ _06585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_143_Left_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10846_ _03686_ _03716_ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13565_ _06510_ _06511_ _06512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10777_ _03572_ _03649_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_54_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12516_ _03556_ net86 net83 _03485_ _05377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13496_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-2\] _06378_ _06437_ _06438_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_82_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12447_ _05301_ _05303_ _05304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_2_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12378_ _05222_ _05228_ _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_1_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07956__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11329_ _04170_ _04171_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10960__B1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12701__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06870_ _05431_ _05452_ _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08381__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13257__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06931__A2 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08540_ _01361_ _01362_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_124_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08471_ _01294_ _01295_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07422_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-20\] _00440_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_106_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07353_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-2\] _00393_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XANTENNA__09633__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10243__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07284_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-1\] _00340_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06998__A2 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09023_ _00394_ _06627_ _06618_ _00398_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_116_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07947__A1 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07947__B2 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09925_ _02731_ _02732_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_141_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10901__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09856_ _02624_ _02739_ _02740_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07175__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08807_ _01628_ _01629_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09787_ _02578_ _02496_ _02575_ _02666_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_06999_ _06059_ _06636_ _06638_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06922__A2 _06081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08738_ _01576_ _01579_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08124__A1 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08124__B2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08669_ _01564_ _01565_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__07214__C _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _03570_ _03573_ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11680_ _00361_ _01610_ _01524_ _00365_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10631_ _03037_ _03430_ _03506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13350_ _06259_ _06262_ _06280_ _06281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_146_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10562_ _03437_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12301_ _05140_ _05144_ _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13281_ _06110_ _06111_ _06109_ _06206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_122_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10493_ net63 _06724_ net57 _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_134_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09388__B1 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12232_ _00354_ _02584_ _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12163_ _05003_ _05004_ _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09157__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11114_ _00384_ _02586_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12094_ _04934_ _04935_ _04937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11045_ _03867_ _03886_ _03887_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08363__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12996_ _05867_ _05896_ _05898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11947_ _04787_ _04788_ _04789_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_98_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08666__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07874__B1 _06523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11878_ net66 net54 _01249_ _01247_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_15_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13617_ _06567_ _06568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10829_ _03572_ _03649_ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11422__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13548_ _00381_ _03727_ _06494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11973__A2 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13479_ _06348_ _06349_ _06420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_112_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07567__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12517__A4 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07929__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ _00871_ _00872_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09710_ _02519_ _02523_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11489__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06922_ _05409_ _06081_ _06103_ _05529_ _06114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12686__B1 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09641_ _02525_ _02526_ _02527_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06853_ _05237_ net170 _05366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10161__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09572_ _00382_ _06679_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08106__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12989__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08523_ _01253_ _01308_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08454_ _01352_ _01307_ _01353_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07405_ _06668_ _00425_ _00426_ _06711_ _05171_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__13890__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08385_ _01285_ _01281_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13402__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07336_ _00380_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_154_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11964__A2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07267_ _05387_ _00324_ _00325_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09006_ _01898_ _01899_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07198_ _06807_ _06808_ _06809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08593__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09908_ _00398_ _00394_ _06674_ _06679_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_09839_ _00376_ _06708_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10152__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12850_ _05728_ _05737_ _05738_ _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11801_ _04614_ _04643_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_96_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12781_ net83 _03725_ _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09845__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11732_ _00378_ _01247_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_139_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13881__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11663_ _04458_ _04459_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XPHY_EDGE_ROW_153_Right_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13402_ _03340_ _00397_ _06336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10614_ _03488_ _03467_ _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11404__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11594_ _04436_ _04185_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_24_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13333_ _06161_ _06166_ _06261_ _06262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_24_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10545_ _03396_ _03403_ _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13157__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07387__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold59_I FreqPhase[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13264_ _03485_ _00384_ _06188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10476_ _03318_ _03319_ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12215_ _00393_ _01610_ _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13195_ _06109_ _06112_ _06113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_90_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12146_ _04966_ _04967_ _04968_ _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07926__A4 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12077_ _04917_ _04918_ _04919_ _04920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11028_ net66 _03266_ _03189_ net54 _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06898__A1 _05811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10694__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12976__B net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12979_ _05876_ _05878_ _05879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08103__A4 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11643__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11643__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13872__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12199__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08170_ _01070_ _01071_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09064__A2 _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11946__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07075__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07121_ _05822_ _06742_ _06743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_119_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07052_ _06624_ _06682_ _06683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07954_ _00851_ _00855_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__12123__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06905_ _05409_ _05919_ _05930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07885_ _00786_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06889__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09624_ _02437_ _02445_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06836_ _05171_ _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XTAP_TAPCELL_ROW_39_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07760__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09555_ _06654_ _06659_ _00398_ _00394_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09827__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08506_ _01402_ _01405_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07838__B1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09486_ _02371_ _02374_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13863__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08437_ _01213_ _01238_ _01335_ _01336_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_92_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08368_ _06618_ _00376_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11937__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07066__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07319_ _00365_ net61 _05182_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08299_ _00935_ _00936_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10330_ _00398_ _00394_ _06701_ _06708_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_33_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10261_ _03139_ _03140_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12000_ _04838_ _04842_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_108_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10192_ _02977_ _02978_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_72_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13951_ _00282_ net101 clknet_leaf_27_clk net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_12902_ _05708_ _05795_ _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13882_ _00213_ net36 clknet_leaf_60_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07541__A2 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12833_ _05546_ _05617_ _05721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09818__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13614__A2 _06563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11625__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12764_ _05597_ _05612_ _05645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_33_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13854__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11715_ net54 _01794_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12695_ _03485_ _00365_ _05571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11646_ net54 _01956_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 net103 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07057__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11577_ _04416_ _04419_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_52_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13316_ _06159_ _06242_ _06244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_141_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10528_ _03355_ _03358_ _03404_ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_24_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13247_ _06154_ _06169_ _06170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10459_ _03253_ _03256_ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_114_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13178_ _05994_ _06093_ _06094_ _06095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12129_ _04889_ _04891_ _04972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07670_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-6\] DDS_Stage.xPoints_Generator1.RegFrequency\[-6\]
+ _00632_ _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09809__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09809__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09340_ _00459_ _02144_ _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_101_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09271_ _02077_ _02128_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07296__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11092__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08222_ _01102_ _01105_ _01101_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_90_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09037__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11919__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07048__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12041__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08153_ net142 _06308_ _06179_ net92 _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07104_ _06713_ _06688_ _06726_ _06727_ _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__12592__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08084_ _00984_ _00985_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_130_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07035_ _05680_ _06668_ _06669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13541__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07220__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08986_ _01812_ _01861_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07937_ _00742_ _00747_ _00838_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07868_ _00749_ _00762_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07523__A2 _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09607_ _02486_ _02494_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07799_ _00715_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ _02346_ _02424_ _02425_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07503__B _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11083__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09469_ _06654_ net58 net95 _06724_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_93_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11500_ _04289_ _04342_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_81_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12480_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-16\] _05338_ _05340_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11431_ _04247_ _04248_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_22_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07039__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12032__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11362_ _04201_ _04202_ _04204_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_61_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13101_ _05852_ _06010_ _06011_ _06012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_21_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10313_ _03112_ _03153_ _03192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11293_ _04133_ _04134_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13032_ _05858_ _05859_ _05857_ _05936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10244_ _02704_ _03122_ _03123_ _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09200__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07211__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10175_ _00373_ _06742_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_89_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13934_ _00265_ net101 clknet_leaf_19_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13865_ _00196_ net36 clknet_leaf_2_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_9_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12816_ _02938_ _00390_ _05703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13796_ _00127_ net36 clknet_leaf_52_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_9_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07278__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12747_ _05533_ _05624_ _05628_ _05629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12678_ _05551_ _05552_ _05553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11629_ _04467_ _04471_ _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_116_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08778__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07575__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12326__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08840_ _01721_ _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07202__A1 _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07202__B2 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08950__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08771_ net137 _06679_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07722_ net108 DDS_Stage.xPoints_Generator1.RegF\[-7\] _00667_ _00676_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11837__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07653_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-8\] _00622_ _00395_ _00623_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07584_ _00566_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09323_ net137 _06710_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07269__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11065__A2 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _01976_ _02056_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08205_ _01102_ _01105_ _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclone39 net139 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_133_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09185_ _02013_ _02041_ _02076_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08136_ _00988_ _01036_ _01037_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07816__I0 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11773__B1 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07441__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08067_ _00967_ _00968_ _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07992__A2 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07018_ _05822_ _06654_ _06655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10328__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08969_ _01706_ _01769_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11980_ _00351_ _02940_ _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10931_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-6\] _03782_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13650_ _06585_ _06591_ _06602_ _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10862_ _03401_ _03707_ _03732_ _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_27_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09249__A2 _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13809__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12601_ _05384_ _05389_ _05468_ _05469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13581_ _06527_ _06528_ _06529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11056__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10793_ _03661_ _03665_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12532_ _04005_ _05392_ _05393_ _05394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_12463_ _04943_ _05320_ _05321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11414_ net66 _02238_ _02236_ net54 _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_50_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12556__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12394_ _05130_ _05163_ _05167_ _05189_ _05246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11345_ _00378_ _01524_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07432__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08775__A4 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11276_ _04116_ _04117_ _04118_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_39_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13015_ _05913_ _05917_ _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10227_ _03106_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_120_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07408__B _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08932__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ _03032_ _03038_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11819__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10089_ _02950_ _02970_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_13917_ _00248_ net36 clknet_3_4__leaf_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_89_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07499__A1 _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13848_ _00179_ net36 clknet_leaf_74_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_58_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13779_ _00114_ clknet_leaf_5_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09660__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09785__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10558__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07423__A1 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09941_ _02718_ _02823_ _02824_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09872_ _02659_ _02665_ _02756_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_5_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07187__B1 _06799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12180__B1 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08923__A1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08823_ _01659_ _01662_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08754_ _01642_ _01650_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07705_ _00666_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__11286__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08685_ _01494_ _01499_ _01582_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07636_ _00606_ _00607_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07567_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[17\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-14\]
+ _00395_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09306_ _02113_ _02114_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12786__A2 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07498_ _05658_ _05724_ _06761_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_36_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ _02077_ _02128_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_62_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12538__A2 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09168_ _01969_ _02057_ _02058_ _02059_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_32_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09403__A2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08119_ net137 _06598_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07414__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11210__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09099_ _01911_ net160 _01991_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_102_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11130_ _00397_ _02238_ _03964_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_101_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XDDS_Module_46 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_11061_ net66 net54 _03340_ _03266_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10012_ _02893_ _02894_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08914__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11963_ net66 _02854_ _02762_ net83 _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08142__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11816__A4 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13702_ _00037_ clknet_leaf_42_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10914_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-14\] _03773_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_82_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11894_ _04519_ _04612_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_129_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10845_ _03686_ _03716_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13633_ _06553_ _06582_ _06583_ _06584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11029__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10776_ _03642_ _03648_ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_hold89_I FreqPhase[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13564_ _06452_ _06509_ _06511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_81_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12515_ _03993_ _03997_ _05375_ _05376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13495_ _06381_ _06436_ _06437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12446_ _04740_ _04741_ _05208_ _05207_ _05205_ _05303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_151_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_97_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07405__A1 _06668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12377_ _05223_ _05227_ _05228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_10_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07956__A2 _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11328_ _04074_ _04098_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10960__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10960__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11259_ _04100_ _04101_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__12701__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10712__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08381__A2 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_74_clk clknet_3_0__leaf_clk clknet_leaf_74_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ _01294_ _01295_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07421_ _06059_ _00438_ _00439_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__A1 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07352_ _00392_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09633__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10243__A3 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07283_ _05182_ _00337_ _00338_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_31_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09022_ _01845_ _01914_ _01915_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09397__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07947__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10951__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ _02804_ _02807_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09855_ _02627_ _02641_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10703__A1 _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08806_ _01625_ _01626_ _01624_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06998_ _05822_ _06637_ _06638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09786_ _02671_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12456__A1 _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08737_ _01560_ _01568_ _01633_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_64_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_65_clk clknet_3_1__leaf_clk clknet_leaf_65_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08124__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08668_ _00385_ _06618_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07619_ _00593_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08599_ _06664_ _00355_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10630_ _03437_ _03501_ _03504_ _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_37_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10561_ _00398_ _00394_ _06724_ _06730_ _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12300_ _05143_ _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_13280_ _06110_ _06111_ _06109_ _06205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10492_ net63 _06724_ net57 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12231_ _04363_ _05072_ _05073_ _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_79_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09388__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09388__B2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11195__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12162_ _05003_ _05004_ _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_20_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11113_ _00387_ net135 _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_92_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12093_ _04934_ _04935_ _04936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_92_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_17_clk_I clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07673__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11044_ _03868_ _03869_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12695__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08363__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07405__C _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12995_ _05881_ _05895_ _05896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_56_clk clknet_3_3__leaf_clk clknet_leaf_56_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11946_ _00393_ _01956_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07874__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__B2 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11877_ net70 _01430_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13616_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-1\] _06508_ _06567_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10828_ _03642_ _03645_ _03647_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_28_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13547_ _00384_ _03725_ _06493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11422__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10759_ _03630_ _03631_ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13478_ _06348_ _06349_ _06419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_42_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09379__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12429_ _05191_ _05209_ _05284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_51_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07929__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07970_ _00823_ _00826_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07583__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06921_ _05409_ _06092_ _05995_ _06103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12686__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11489__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12686__B2 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10697__B1 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09640_ net138 _06742_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06852_ _05291_ _05313_ _05335_ net129 _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_93_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09571_ _02379_ _02457_ _02458_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08106__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_47_clk clknet_3_4__leaf_clk clknet_leaf_47_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08522_ _01351_ _01421_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__12989__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08453_ _01255_ _01300_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_147_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07404_ _06668_ _06693_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08384_ _01282_ _01283_ _01284_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_129_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07335_ _00378_ _00379_ _05182_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12610__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11964__A3 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ _05182_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-4\] _00325_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09005_ _06659_ _00376_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07197_ _06726_ _06759_ _06774_ _06703_ _06146_ _06808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_130_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11177__A1 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08593__A2 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09790__A1 _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09907_ _00398_ _06674_ _06679_ _00394_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12677__A1 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ _00379_ _06701_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10152__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09769_ _02509_ _02570_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11800_ _04623_ _04641_ _04642_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12780_ _05659_ _05568_ _05566_ _05663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09845__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11731_ _04572_ _04573_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11662_ _04484_ _04503_ _04504_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_95_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13401_ _06244_ _06251_ _06334_ _06335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10613_ _03419_ _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_12_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11593_ _00390_ _01247_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11404__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10544_ _03360_ _03395_ _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13332_ _06158_ _06260_ _06261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13157__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10475_ _03344_ _03351_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13263_ net147 _00387_ _06187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12214_ _00390_ _01693_ _05057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08033__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13194_ _06110_ _06111_ _06112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10915__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12145_ _04965_ _04973_ _04988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12076_ net86 net83 _02762_ _02586_ _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__12668__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11027_ _03867_ _03868_ _03869_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_108_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11340__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07544__B1 _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_29_clk clknet_3_7__leaf_clk clknet_leaf_29_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_91_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12976__C _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12978_ _05764_ _05877_ _05878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11643__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11929_ _00378_ _02238_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12199__A3 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07120_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[4\] _06742_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_125_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07075__A2 _06700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07051_ _05583_ _06681_ _06682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10906__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07953_ _00852_ _00853_ _00854_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_128_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06904_ _05897_ _05908_ _05919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07884_ _06637_ net58 _00355_ _06633_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09623_ _02437_ _02445_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06835_ net1 _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XTAP_TAPCELL_ROW_39_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06889__A2 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone56_I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09554_ _06654_ _00398_ _00394_ _06659_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09827__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08505_ _01403_ _01404_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07838__A1 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07838__B2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09485_ _02372_ _02373_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_53_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08436_ _01143_ _01096_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_18_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08367_ _06598_ _00379_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11398__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07318_ _00366_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XANTENNA__11937__A3 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08298_ _01182_ _01183_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07249_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-7\] _00310_ _05182_ _00311_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10260_ _00376_ _06742_ _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10191_ _03027_ _03071_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_72_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13950_ _00281_ net101 clknet_leaf_26_clk net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07236__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12901_ _05712_ _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13881_ _00212_ net36 clknet_leaf_62_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_12832_ _05641_ _05643_ _05719_ _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_17_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09818__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07829__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12822__A1 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11625__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12763_ _05597_ _05612_ _05644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_84_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11714_ net66 _01956_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12694_ net148 _00369_ _05570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11645_ _04485_ _04486_ _04487_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11389__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 net107 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11576_ _04417_ _04418_ _04176_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_25_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13315_ _00369_ _03727_ _06060_ _06242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10527_ _03396_ _03403_ _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_134_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13246_ _06158_ _06167_ _06169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10458_ _00522_ _03328_ _03335_ _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_123_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13177_ _05996_ _05997_ _06094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10389_ _03263_ _03265_ _03267_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11561__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12128_ _04966_ _04969_ _04970_ _04971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13790__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12059_ _04899_ _04900_ _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09809__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09270_ _02073_ _02074_ _02160_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08221_ _01098_ _01122_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13369__A2 _06208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08152_ _01052_ _01053_ _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07048__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12041__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07103_ _05420_ _05485_ _06232_ _06727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08083_ _06179_ _00370_ _00982_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_9_clk clknet_3_3__leaf_clk clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07034_ _05647_ _05409_ _06668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_141_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13541__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11552__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_149_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08985_ _01812_ _01861_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07936_ _00737_ _00748_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07867_ _00764_ _00765_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09606_ _02489_ _02493_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07798_ net58 DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[16\] _00395_ _00715_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09537_ net61 net142 _06701_ _06708_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__07503__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08484__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09468_ _06654_ net95 _06724_ net58 _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_109_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08419_ _01319_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09399_ _02286_ _02287_ _02288_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_124_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11430_ _04204_ _04271_ _04272_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08236__A1 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07039__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12032__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11361_ _04203_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13100_ _05854_ _06009_ _06011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_105_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10312_ _03082_ _03162_ _03160_ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11292_ _04133_ _04134_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_120_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10243_ net63 _06701_ net57 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_13031_ _05822_ _05934_ _05935_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10174_ _03053_ _03054_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06970__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07681__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13933_ _00264_ net101 clknet_leaf_14_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_88_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13864_ _00195_ net36 clknet_leaf_63_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_44_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12815_ _02854_ _00393_ _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13795_ _00126_ net36 clknet_leaf_66_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_56_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08475__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12746_ _05530_ _05532_ _05628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12677_ net135 _00397_ _05512_ _05552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_71_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11628_ _04468_ _04470_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10034__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08778__A2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11559_ _00397_ _01249_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11782__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13229_ _05959_ _06061_ _05953_ _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08950__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08770_ _00355_ _06674_ _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13287__A1 _06131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06961__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07721_ _00675_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11837__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13039__A1 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ DDS_Stage.xPoints_Generator1.CosNew\[-8\] _00621_ _00577_ _00622_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07583_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[25\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-6\]
+ _00395_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _00355_ _06708_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07269__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09253_ _00459_ _02144_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_35_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone18 net90 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08204_ _01102_ _01105_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09184_ _02016_ _02040_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08135_ _01018_ _01035_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11773__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07766__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11773__B2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08066_ _00771_ _00799_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07441__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07017_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-11\] _06654_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11525__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08968_ _01801_ _01803_ _01862_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__06952__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07919_ _00801_ _00819_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08899_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[7\] _01794_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_3_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10930_ _03781_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10861_ _03730_ _03731_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12600_ _05379_ _05383_ _05468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13580_ _06237_ _06239_ _06476_ _06528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_10792_ _03082_ _03664_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_38_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12531_ _04006_ _04007_ _05393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12462_ _05016_ _05316_ _05238_ _05320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11413_ _04245_ _04249_ _04255_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12393_ _05130_ _05163_ _05245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11344_ _04180_ _04184_ _04186_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_132_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11275_ _00393_ _02051_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11516__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_148_Right_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13014_ _05914_ _05915_ _05916_ _05917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_10226_ _03080_ _03082_ _03078_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13745__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ _03034_ _03037_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08932__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09904__B _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06943__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11819__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10088_ _02961_ _02969_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13916_ _00247_ net36 clknet_leaf_42_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_57_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_126_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13847_ _00178_ clknet_leaf_42_clk DDS_Stage.xPoints_Generator1.RegP\[-1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13778_ _00113_ clknet_leaf_15_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12729_ _03018_ _00381_ _05609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12492__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10558__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08620__A1 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07423__A2 _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09940_ _02721_ _02735_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_110_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09871_ _02654_ _02658_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_110_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13736__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12180__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12180__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08822_ _01642_ _01650_ _01717_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08923__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06934__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08753_ _01645_ _01649_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_135_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07704_ net36 _05237_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08684_ _01489_ _01493_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08687__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10494__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07635_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-11\] DDS_Stage.xPoints_Generator1.RegFrequency\[-11\]
+ _00602_ _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07566_ _00557_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10246__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09305_ _02113_ _02114_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_35_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07497_ _06146_ _05745_ _00501_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_119_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09236_ _02098_ _02127_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09167_ _01976_ _02056_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_16_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09403__A3 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08118_ _01006_ _01014_ _01019_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09098_ _01913_ _01937_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08049_ _00949_ _00950_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11060_ net66 _03340_ _03266_ net54 _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_102_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDDS_Module_47 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__07178__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13727__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10011_ _02712_ _02794_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08914__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_48_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11962_ _00359_ _02586_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13701_ _00036_ clknet_leaf_53_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__A3 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10913_ _05822_ _06811_ _03772_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11893_ _04520_ _04613_ _04733_ _04735_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_86_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13632_ _06526_ _06552_ _06583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10844_ _03688_ _03690_ _03715_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_128_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11029__A3 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10237__A1 _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13563_ _06452_ _06509_ _06510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10775_ _03645_ _03647_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07102__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12514_ _03988_ _03992_ _05375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_57_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__A1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13494_ _06314_ _06435_ _06436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12445_ _05202_ _05203_ _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12376_ _05063_ _05067_ _05224_ _05225_ _05227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_2_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07956__A3 _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11327_ _04146_ _04168_ _04169_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__10960__A2 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11258_ _03852_ _03969_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07169__A1 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10209_ _03085_ _03089_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11189_ _04015_ _04017_ _04031_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_82_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13662__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07420_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-21\] _00439_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13414__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07892__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07351_ _00390_ net63 _05182_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07282_ _06081_ _06788_ _06146_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09021_ net138 net96 _06627_ _06691_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_26_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09397__A2 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13957__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10400__A1 _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10951__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09923_ _02805_ _02806_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_84_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09854_ _02627_ _02641_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06907__A1 _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11900__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08805_ net56 _01348_ _01700_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09785_ _02586_ _02670_ _00395_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06997_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-14\] _06637_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08736_ _01563_ _01567_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10467__A1 _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08667_ _00388_ _06598_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07618_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\] _00592_ _00395_ _00593_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_64_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08598_ _01495_ _01496_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_93_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10219__A1 _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07549_ _05182_ _00542_ _00544_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__11967__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10560_ _00398_ _06724_ _06730_ _00394_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09219_ _02030_ _02038_ _02110_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10491_ _03364_ _03367_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11719__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12230_ net87 net84 _02584_ _02499_ _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09388__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13948__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07399__A1 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11195__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12161_ _04915_ _04928_ _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07239__B _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11112_ _03838_ _03953_ _03954_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_92_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12092_ _04802_ _04844_ _04935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_11043_ _03868_ _03869_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12695__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12994_ _05884_ _05894_ _05895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11945_ _00390_ _02051_ _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__A2 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11876_ _04704_ _04718_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13615_ _06516_ _06564_ _06565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10827_ _03697_ _03698_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13546_ _06423_ _06489_ _06490_ _06492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10758_ _03596_ _03601_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13477_ _06417_ _06418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_124_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10689_ _03561_ _03562_ _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12428_ _05223_ _05227_ _05283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09379__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13939__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12359_ _05205_ _05207_ _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_11_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06920_ _05431_ _05463_ _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__12686__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10697__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10697__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06851_ _05182_ _05302_ net17 _05204_ _05346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_93_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07562__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09570_ _02380_ _02381_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_117_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13635__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08106__A3 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08521_ _01354_ _01420_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08452_ _01255_ _01300_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_46_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07403_ _05529_ _06666_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_9_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08383_ _06642_ _00363_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07334_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-7\] _00379_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_128_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12610__A2 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07265_ _00321_ _00323_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11964__A4 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09004_ _06654_ _00379_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07196_ _05702_ _06806_ _05658_ _05669_ _06807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_115_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11177__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07774__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09790__A2 _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09906_ _02788_ _02704_ _02789_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_74_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12677__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ _00373_ _06710_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07553__A1 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09768_ _02589_ _02653_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08719_ _01537_ _01601_ _01615_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_69_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09699_ _02581_ _02583_ _02585_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xrebuffer60 _00366_ net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11730_ _04492_ _04494_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06917__I _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11661_ _04501_ _04502_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07241__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13400_ _06241_ _06252_ _06334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10612_ _03422_ _03466_ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07608__A2 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11592_ _04425_ _04433_ _04434_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13331_ _06167_ _06260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10543_ _03082_ _03402_ _03418_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13262_ _06096_ _06184_ _06185_ _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_94_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10474_ _03345_ _03342_ _03350_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12213_ _00397_ _01524_ _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08033__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13193_ _05936_ _06007_ _06111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12144_ _04959_ _04977_ _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_103_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12117__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12075_ net86 _02762_ _02586_ net83 _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_21_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11026_ _00361_ _03018_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07544__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11340__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12977_ net70 _03727_ _05877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09297__A1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11928_ _04766_ _04769_ _04770_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11859_ _04694_ _04695_ _04701_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12199__A4 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13529_ _06239_ _06404_ _06237_ _06473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07050_ _06232_ _05485_ _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_125_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_63_clk_I clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09221__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07952_ net143 _06633_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_78_clk_I clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06903_ _05572_ _05463_ _05908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07883_ _00774_ _00783_ _00784_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07535__A1 _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ _02507_ _02508_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06834_ _05139_ DDS_Stage.LCU.state\[0\] _05160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13608__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09553_ _02351_ _02439_ _02440_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09288__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09827__A3 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08504_ net137 _06664_ net95 _06308_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11095__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07838__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09484_ _00376_ _06685_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08435_ _01236_ _01165_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_77_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_16_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ _06627_ _00373_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11398__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07317_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-11\] _00366_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_34_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08297_ _01179_ _01191_ _01198_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_2_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11937__A4 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_12_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07248_ _05658_ _00307_ _00308_ _00309_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_143_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _05182_ _06791_ _06792_ _06793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__10923__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10190_ _03049_ _03070_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07526__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12900_ _05757_ _05793_ _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_21_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13880_ _00211_ net36 clknet_leaf_61_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_12831_ _05651_ _05718_ _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_97_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12762_ _05554_ _05615_ _05642_ _05643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07829__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12822__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11713_ _04547_ _04554_ _04555_ _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12693_ _05564_ _05565_ _05568_ _05569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_84_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11644_ net66 net54 _01956_ _01794_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_65_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11389__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11575_ _00384_ _01249_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_30_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput16 net105 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13314_ _06163_ _06164_ _06240_ _06241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10526_ _03082_ _03402_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13245_ _06161_ _06166_ _06167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10457_ _03182_ _03330_ _03334_ _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_0_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13176_ _05996_ _05997_ _06093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10388_ _05280_ _03266_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11561__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12127_ _04967_ _04968_ _04970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12058_ _04899_ _04900_ _04901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11009_ _03849_ _03851_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10824__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08220_ _01111_ _01112_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08151_ _01050_ _01051_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09442__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07102_ _05572_ _05431_ _06726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_113_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08082_ _06179_ _00370_ _00982_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_99_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07033_ _05897_ _06666_ _06667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13887__CLK clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11552__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08984_ _01876_ _01877_ _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_149_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07935_ _00827_ _00836_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07508__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone8_I net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07866_ _00767_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_138_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09605_ _02318_ _02392_ _02490_ _02491_ _02492_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_3_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07797_ _00714_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09536_ net61 _06701_ _06708_ net142 _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10815__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09467_ _02342_ _02355_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_109_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08484__A2 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09681__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08418_ _01249_ _01318_ _00395_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09398_ net58 _06724_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08349_ _00870_ _00873_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_46_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08236__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12032__A3 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11240__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11360_ _00378_ _01610_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10311_ _05822_ _03188_ _03190_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11291_ _04053_ _04055_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_132_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13030_ _05280_ net32 _05935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10242_ net63 _06701_ net57 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08944__B1 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10173_ _02885_ _02968_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07211__A3 _06787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13932_ _00263_ net101 clknet_leaf_19_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_13863_ _00194_ net36 clknet_leaf_64_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_0_88_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12814_ _02762_ _00397_ _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13794_ _00125_ net36 clknet_leaf_65_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_85_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12745_ _05438_ _05624_ _05625_ _05626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_139_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08475__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12676_ _05510_ _05511_ _05551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_127_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ _04467_ _04469_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_41_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10034__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11558_ _04396_ _04400_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_123_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11782__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10509_ _03303_ _03304_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_122_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11489_ _00387_ _01524_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13228_ _06147_ _06148_ _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13159_ _06071_ _06072_ _06073_ _06074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_85_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06961__A2 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07720_ net104 DDS_Stage.xPoints_Generator1.RegF\[-8\] _00667_ _00675_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07651_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-8\] DDS_Stage.xPoints_Generator1.RegFrequency\[-8\]
+ _00620_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13039__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07910__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07582_ _00565_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12798__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09321_ _02207_ _02211_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_146_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09252_ _02139_ _02143_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_8_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08203_ _01103_ _01104_ _00993_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_16_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09183_ _02073_ _02074_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08134_ _01018_ _01035_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_71_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11773__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08065_ _00951_ _00965_ _00966_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_56_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07441__A3 _06125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07016_ _06146_ _06652_ _06653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11525__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07782__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08967_ _01810_ _01812_ _01861_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_07918_ _00801_ _00819_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08898_ _06059_ _01791_ _01793_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08154__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07849_ _06308_ _00376_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10860_ _03654_ _03703_ _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09519_ _05182_ _02407_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10791_ _03401_ _03663_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_149_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12530_ _04006_ _04007_ _05392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11461__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06925__I _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12461_ _05293_ _05315_ _05318_ _05319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09406__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11412_ _04240_ _04244_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12392_ _05164_ _05190_ _05242_ _05243_ _05244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_151_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12961__A1 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11343_ _00390_ _01247_ _04185_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_104_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11274_ _00390_ _02153_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13013_ _03340_ _00381_ _05916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11516__A2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10225_ _03019_ _03105_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08393__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_3__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _03036_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_100_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06943__A2 _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10087_ _02885_ _02968_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13915_ _00246_ net36 clknet_leaf_53_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_89_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_113_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09893__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12229__B1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13846_ _00177_ clknet_leaf_42_clk DDS_Stage.xPoints_Generator1.RegP\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13777_ _00112_ clknet_leaf_20_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10989_ _03829_ _03830_ _03831_ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__11452__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12728_ _02940_ _00384_ _05608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12659_ _05434_ _05437_ _05533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11204__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10558__A3 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08620__A2 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09870_ _02754_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_5_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12180__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ _01645_ _01649_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06934__A2 _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08752_ _01646_ _01647_ _01648_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_07703_ _00665_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08683_ _01481_ _01580_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08687__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07634_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-11\] DDS_Stage.xPoints_Generator1.RegFrequency\[-11\]
+ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07565_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[16\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-15\]
+ _00395_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_24_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clone31_I net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09304_ _02106_ _02107_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10246__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07496_ _06232_ _06713_ _05897_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_146_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _02101_ _02126_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09166_ _01972_ _01947_ _01971_ _02047_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__06870__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08117_ _01009_ _01013_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09403__A4 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09097_ _01988_ _01989_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10954__B1 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08048_ _00355_ _06618_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDDS_Module_37 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__07178__A2 _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDDS_Module_48 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10010_ _02790_ _02793_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09999_ net63 _06685_ _02608_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08127__A1 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11961_ _04766_ _04767_ _04768_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09875__A1 _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13700_ _00035_ clknet_leaf_64_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10912_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-15\] _03772_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08142__A4 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11892_ _04730_ _04731_ _04734_ _04611_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_13631_ _06560_ _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_129_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10843_ _03696_ _03714_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11029__A4 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11434__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13562_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-1\] _06508_ _06509_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10774_ _00398_ _06742_ _03646_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_55_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07102__A2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12513_ _03999_ _04010_ _05373_ _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_13493_ _06385_ _06434_ _06435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08850__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07687__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12444_ _05298_ _05208_ _05299_ _05300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12375_ _05119_ _05129_ _05225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_10_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11326_ _04166_ _04167_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_120_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07956__A4 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11257_ _04074_ _04098_ _04099_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08366__A1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07169__A2 _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10208_ _03087_ _03088_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_11188_ _04022_ _04030_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_128_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10139_ _02995_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_141_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13662__A2 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13829_ _00160_ clknet_leaf_48_clk DDS_Stage.xPoints_Generator1.RegF\[-4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13414__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07350_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-3\] _00391_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07170__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07281_ _05658_ _06624_ _00336_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_116_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09020_ net96 _06627_ _06691_ net138 _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_139_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_152_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09922_ _00376_ _06710_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09554__B1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ _02690_ _02737_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11900__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08804_ _01425_ _01507_ _01605_ _01687_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_147_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09784_ _02666_ _02669_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08109__A1 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06996_ _06146_ _06635_ _06636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08735_ _01571_ _01598_ _01631_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09857__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08666_ _06627_ _00382_ _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07617_ DDS_Stage.xPoints_Generator1.CosNew\[-13\] _00591_ _00577_ _00592_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_81_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13893__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08597_ net97 net153 _06672_ net137 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_37_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07548_ _05658_ _06661_ _00543_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_76_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11967__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07096__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07479_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-11\] _00487_ _00488_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09218_ _02033_ _02037_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10490_ _03037_ _03366_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_134_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07300__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12916__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11719__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ _02013_ _02041_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_121_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08596__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12160_ _04988_ _05001_ _05002_ _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11111_ _03839_ _03840_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12091_ _04914_ _04932_ _04933_ _04934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_92_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11042_ _03829_ _03883_ _03884_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07020__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12993_ _05893_ _05894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11944_ _00397_ _01794_ _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13884__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11875_ _04717_ _04703_ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10826_ _03652_ _03659_ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13614_ _06519_ _06563_ _06564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07087__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10757_ _03565_ _03595_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13545_ _06424_ _06425_ _06490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_138_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13476_ _06412_ _06415_ _06417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_153_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10688_ _03529_ _03534_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12907__A1 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12427_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-15\] _05281_ _05282_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_106_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13580__A1 _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12358_ _04224_ _04412_ _05206_ _05207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_22_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11309_ _04149_ _04150_ _04151_ _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12289_ _04396_ _05131_ _05132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09536__B1 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06850_ _05324_ _05291_ _05335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10697__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09839__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13635__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08520_ _01363_ _01419_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11646__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08106__A4 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08511__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13875__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08451_ _01303_ _01305_ _01350_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_148_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07402_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-24\] _00424_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_46_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08382_ _00367_ _06637_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07078__A1 _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07333_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-7\] _00378_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_144_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08814__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07264_ _05658_ _06826_ _00322_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_27_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09003_ _06664_ _00373_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07195_ _05409_ _05452_ _06806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_130_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09905_ net63 _06679_ _02608_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_74_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11334__B1 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09836_ _02719_ _02720_ _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07790__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08750__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07553__A2 _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06979_ _05420_ _05431_ _06621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09767_ _02591_ _02644_ _02652_ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_69_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08718_ _01540_ _01600_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07803__B _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09698_ _05280_ net135 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer50 _02610_ net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_83_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08502__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer61 _01938_ net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13866__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08649_ _06649_ _00370_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11660_ _04501_ _04502_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07069__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10611_ _05822_ _03484_ _03486_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11591_ _04431_ _04432_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08805__A2 _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13330_ _06183_ _06192_ _06258_ _06259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10542_ _03399_ _03401_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06933__I _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13261_ _06097_ _06098_ _06185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_94_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10473_ _03259_ _03260_ _03346_ _03348_ _03349_ _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_33_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08569__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12212_ _05051_ _05054_ _05055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13192_ _05938_ _06005_ _06110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12143_ _04979_ _04982_ _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07241__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12117__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12074_ _00359_ _02584_ _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11025_ _00365_ _02940_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08741__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12976_ _05765_ _05874_ net70 _03727_ _05876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_87_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13857__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11927_ _04767_ _04768_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_59_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11858_ _04676_ _04690_ _04691_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_129_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10809_ _03668_ _03669_ _03667_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_31_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12053__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11789_ _04628_ _04631_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_28_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13528_ _06407_ _06431_ _06471_ _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13459_ _06397_ _06398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07232__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07951_ net74 _06627_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06902_ _05420_ _05886_ _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07882_ net157 _00782_ _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11867__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08732__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06833_ _05139_ DDS_Stage.LCU.state\[0\] DDS_Stage.LCU.state\[1\] DDS_Stage.LCU.SelMuxConfig
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09621_ _02469_ _02476_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13608__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09552_ _02352_ _02353_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09288__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08503_ net58 _06664_ net95 _06308_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__09827__A4 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13848__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08496__B1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ _00379_ _06679_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11095__A2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08434_ _01332_ _01333_ _01236_ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08365_ _01263_ _01264_ _01265_ _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_92_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_rebuffer41_I net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07316_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-11\] _00365_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
XFILLER_0_117_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08296_ _01181_ _01190_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07471__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07247_ _05409_ _06447_ _06733_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_117_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _06146_ _05886_ _06645_ _06629_ _06792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_42_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07223__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11307__B1 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09819_ _02703_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_12830_ _05654_ _05717_ _05718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07252__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12761_ _05556_ _05614_ _05642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11712_ net66 net54 _01794_ _01792_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_12692_ _05566_ _05567_ _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_139_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12035__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11643_ net66 _01956_ _01794_ net54 _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09987__B1 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11574_ _00381_ _01430_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 net128 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10525_ _03399_ _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13313_ _00378_ _03558_ _06165_ _06240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_24_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07462__A1 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07695__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13244_ _06162_ _06165_ _06166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_hold57_I FreqPhase[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10456_ _03333_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13175_ _06087_ _06090_ _06091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07214__B2 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[23\] _03266_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12126_ _04967_ _04968_ _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07427__C _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12057_ _04761_ _04763_ _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08714__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07517__A2 _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11008_ _03792_ _03794_ _03848_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_88_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12959_ _05797_ _05855_ _05856_ _05857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_48_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08150_ _01050_ _01051_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10588__A1 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09442__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07101_ _06059_ _06723_ _06725_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08081_ _06179_ _00370_ _00982_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_43_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07453__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07032_ _05572_ _05669_ _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07205__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11552__A3 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08983_ _06664_ _00370_ _01808_ _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_149_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07934_ _00830_ _00835_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07508__A2 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07865_ _00736_ _00763_ _00766_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10512__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09604_ _02391_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_155_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07796_ DDS_Stage.xPoints_Generator1.RegFrequency\[-1\] DDS_Stage.xPoints_Generator1.RegF\[-1\]
+ _00402_ _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09535_ _02350_ _02354_ _02422_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09466_ _02350_ _02354_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_148_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09681__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ _00418_ _01317_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09397_ _06654_ net96 _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08348_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[1\] _01249_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_117_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12032__A4 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07444__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08279_ _01083_ _01091_ _01180_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11240__A2 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10310_ _05280_ _03189_ _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11290_ _04128_ _04131_ _04132_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10241_ _03117_ _03120_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_30_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08944__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10172_ _02964_ _02967_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08944__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13931_ _00262_ net101 clknet_leaf_19_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_88_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13862_ _00193_ net36 clknet_leaf_42_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_12813_ _05697_ _05698_ _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13793_ _00124_ net36 clknet_leaf_66_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_clkbuf_leaf_62_clk_I clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12744_ _05530_ _05532_ _05625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12675_ _05505_ _05547_ _05548_ _05549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11626_ _00372_ _01524_ _01430_ _00375_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_154_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_77_clk_I clknet_3_2__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07435__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11557_ _04397_ _04398_ _04399_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__13508__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10508_ _03303_ _03304_ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11488_ _00381_ _01693_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13227_ _06063_ _06077_ _06148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10439_ _03221_ _03236_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13158_ _00372_ _03679_ _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12109_ _04873_ _04951_ _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13089_ _05993_ _05998_ _05999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_15_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10799__B _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09360__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07650_ _00618_ _00619_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_144_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07910__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07581_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[24\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-7\]
+ _00395_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09320_ _02208_ _02209_ _02210_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__12798__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09251_ _02140_ _02141_ _02142_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_118_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08202_ net91 _05398_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09182_ _00370_ _06679_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08133_ _01005_ _01020_ _01034_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_44_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07426__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08064_ _00963_ net72 _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07015_ _06651_ _06629_ _06652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09179__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08966_ _01832_ _01860_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07917_ _00788_ _00818_ _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08897_ _05280_ _01792_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08154__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07848_ net152 _00373_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclone2 net62 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XANTENNA__12238__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10929__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07779_ _00705_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_27_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09518_ _02395_ _02405_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10790_ _03586_ _03593_ _03662_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11461__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ _02273_ _02301_ _02337_ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12460_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-19\] _05317_ _05290_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-20\]
+ _05318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_53_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09406__A2 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11411_ _04251_ _04252_ _04253_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07417__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12391_ _05192_ _05201_ _05205_ _05207_ _05243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_62_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11342_ _04180_ _04184_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12961__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11273_ _00397_ _01956_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13012_ _03266_ _00384_ _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11516__A3 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10224_ _05387_ _03103_ _03104_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_101_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08393__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10155_ _02779_ _03035_ _03031_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_7_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10086_ _02964_ _02967_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12477__A1 _05336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13727__CLK clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13914_ _00245_ net36 clknet_leaf_53_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_96_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09893__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12229__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13845_ _00176_ clknet_leaf_45_clk DDS_Stage.xPoints_Generator1.RegP\[-3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12229__B2 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13776_ _00111_ clknet_leaf_22_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10988_ _00375_ _02762_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12727_ _02938_ _00387_ _05607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11452__A2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12658_ _03977_ _05433_ _05531_ _05532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_37_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07408__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11609_ _04442_ _04450_ _04451_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11204__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12589_ _05411_ _05426_ _05456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_10_clk clknet_3_3__leaf_clk clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08081__A1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07168__B _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08820_ _01653_ _01681_ _01715_ _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_146_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08751_ _06627_ _00385_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77_clk clknet_3_2__leaf_clk clknet_leaf_77_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07702_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-1\] _00664_ _00395_ _00665_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08682_ _01579_ _01576_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07633_ _00605_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07564_ _00556_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09303_ _02109_ _02125_ _02193_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10246__A3 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07495_ _00500_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09234_ _02109_ _02125_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_145_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09165_ _01976_ _02056_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13196__A2 _05840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06870__A2 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08116_ _00989_ _01016_ _01017_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12943__A2 _05840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09096_ _00370_ _06674_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10954__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10954__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08047_ net138 _06627_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10706__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDDS_Module_38 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XDDS_Module_49 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_101_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07178__A3 _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ net63 _06685_ _02608_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08949_ _01754_ _01762_ _01843_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08127__A2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_68_clk clknet_3_0__leaf_clk clknet_leaf_68_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09324__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11960_ _04765_ _04777_ _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10911_ _03771_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07886__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11891_ _04600_ _04605_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13630_ _06546_ _06580_ _06581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07541__B _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10842_ _03699_ _03713_ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11434__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13561_ _06454_ _06507_ _06508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10773_ _03644_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_149_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12512_ _03985_ _03998_ _05373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13492_ _06391_ _06433_ _06434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12443_ _04740_ _04741_ _05208_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-25\]
+ _05299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__11198__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12374_ _05119_ _05129_ _05224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10945__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11325_ _04166_ _04167_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_127_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11256_ _04096_ _04097_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08366__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _02943_ _03002_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11187_ _04025_ _04029_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_128_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10138_ _05822_ _03018_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_59_clk clknet_3_3__leaf_clk clknet_leaf_59_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09315__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10069_ _02872_ _02875_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_141_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07877__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12870__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13828_ _00159_ clknet_leaf_49_clk DDS_Stage.xPoints_Generator1.RegF\[-5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_106_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13759_ _00094_ clknet_leaf_78_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07280_ _05734_ _06681_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08054__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09921_ _00379_ _06708_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12689__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09554__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09554__B2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09852_ _02736_ _02716_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08803_ _01695_ _01698_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09783_ _02668_ _02582_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06995_ _05507_ _06221_ _06383_ _06635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08109__A2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08734_ _01574_ _01597_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11113__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09857__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13653__A3 _06605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08665_ _01467_ _01561_ _01562_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06915__I0 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07616_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\] DDS_Stage.xPoints_Generator1.RegFrequency\[-13\]
+ _00590_ _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08596_ net58 net95 net152 _06672_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_48_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_132_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07547_ _05951_ _06704_ _00479_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07788__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07096__A2 _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07478_ _05171_ _00485_ _00486_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_119_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09217_ _02102_ _02105_ _02108_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_17_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12916__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11719__A3 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09148_ _02016_ _02040_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08596__A2 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09079_ _01863_ _01866_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11110_ _03839_ _03840_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12090_ _04930_ _04931_ _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_141_Left_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_92_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11041_ _03830_ _03831_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09545__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11352__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12992_ _05888_ _05892_ _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11943_ _04782_ _04785_ _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_54_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07271__B _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11874_ _04715_ _04716_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_95_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13613_ _06467_ _06562_ _06563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10825_ _03636_ _03651_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13544_ _06424_ _06425_ _06489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_hold87_I FreqPhase[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07087__A2 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10756_ _03401_ _03599_ _03628_ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__I0 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13475_ _06413_ _06414_ _06415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10687_ _03496_ _03528_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12426_ _04174_ _05276_ _05281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12907__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13580__A2 _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12357_ _04345_ _04411_ _05206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11308_ net86 net83 _02940_ _02938_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_120_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12288_ _04400_ _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_120_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09536__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09536__B2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11239_ _00351_ _03189_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11343__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09839__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11646__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12843__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08511__A2 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08450_ _06633_ _00370_ _01306_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_9_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07401_ _05387_ _00418_ _00423_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08381_ _06649_ _00357_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07332_ _00377_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10082__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07263_ _05409_ _05875_ _06666_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09002_ _01835_ _01894_ _01895_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07194_ _06805_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09224__B1 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09904_ net63 _06679_ _02608_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11334__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11334__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09835_ _02535_ _02619_ _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08750__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13087__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09766_ _02650_ _02651_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06978_ _05908_ _06620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08717_ _01613_ _01606_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09697_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[15\] _02584_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xrebuffer40 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-15\] net139 vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xrebuffer51 _02600_ net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__08502__A2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer62 net73 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_08648_ _01542_ _01545_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_95_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08579_ net58 _06664_ net95 _06308_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10937__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10610_ _05280_ _03485_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11590_ _04431_ _04432_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_9_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10073__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10541_ _03414_ _03415_ _03417_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08018__A1 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13260_ _06097_ _06098_ _06184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13011__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10472_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-2\] _03347_ _03349_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_150_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12211_ _04945_ _05053_ _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08569__A2 _06523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13191_ _06041_ _06108_ _06109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12142_ _04984_ _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07241__A2 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12117__A3 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12073_ _04894_ _04895_ _04896_ _04916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10128__A2 _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11024_ _00369_ _02938_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08741__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13078__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12975_ net70 _03725_ _05764_ _05874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11926_ _04767_ _04768_ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11857_ _04644_ _04699_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_74_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10808_ _03676_ _03678_ _03680_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08257__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12053__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09454__B1 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11788_ _04629_ _04630_ _04541_ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__07304__I0 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13527_ _06395_ _06406_ _06471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10739_ _03540_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13458_ _00378_ _03727_ _06324_ _06397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_23_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12409_ _04866_ _05251_ _05262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11013__B1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13389_ _00372_ _00375_ _03727_ _06323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_10_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13793__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09509__A1 _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07950_ _00357_ _06637_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08980__A2 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06991__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ _05431_ _05463_ _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07881_ _00782_ _00778_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11867__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08732__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09620_ _02419_ _02468_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06832_ DDS_Stage.LCU.state\[2\] _05139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09551_ _02352_ _02353_ _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12816__A1 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08502_ _00355_ _06659_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08496__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09482_ _00373_ _06691_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08496__B2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11095__A3 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08433_ _01096_ _01144_ _01238_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_37_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08248__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13241__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08364_ net153 _00385_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07315_ _00364_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08295_ _01195_ _01193_ _01196_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_rebuffer34_I net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07246_ _06232_ _05474_ _05658_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_116_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07471__A2 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07177_ _06787_ _06788_ _05658_ _06790_ _06791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_76_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11555__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13784__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11307__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11307__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06982__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09818_ _00355_ _06744_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09920__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07931__B1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09749_ _02554_ _02633_ _02634_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12760_ _05551_ _05552_ _05549_ _05641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_87_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11711_ net66 _01794_ _01792_ net54 _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_68_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12691_ net54 _03679_ _03725_ net86 _05567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_65_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11642_ net70 _01792_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12035__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09987__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09987__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11573_ _04414_ _04415_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_65_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput18 net124 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13312_ _06237_ _06238_ _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_10524_ _03308_ _03400_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__07462__A2 _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13243_ _06163_ _06164_ _06165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10455_ _03255_ _03331_ _03332_ _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_122_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13174_ _06088_ _06089_ _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10386_ _05182_ _03264_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_131_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12125_ _00365_ _02409_ _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13299__A1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12056_ _04894_ _04897_ _04898_ _04899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11007_ _03849_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12958_ _05801_ _05816_ _05856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11909_ _04748_ _04751_ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12889_ _05671_ _05672_ _05782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_28_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10037__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09978__A1 _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07989__B1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07100_ _05822_ _06724_ _06725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08080_ _05833_ _05398_ _00376_ _00373_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_99_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07031_ _06059_ _06663_ _06665_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11537__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11552__A4 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ _01875_ _01807_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06964__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_71_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07933_ _00831_ _00834_ _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07864_ _00764_ _00765_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10512__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09603_ _02155_ _02225_ _02311_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_79_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07795_ _00713_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clone54_I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09534_ _02345_ _02349_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10276__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09465_ _02351_ _02352_ _02353_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07141__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08416_ _01314_ _01316_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_47_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09396_ _00355_ _06710_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08347_ _01245_ _01246_ _01248_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07796__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08278_ _01085_ _01090_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07444__A2 _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07229_ _06714_ _06666_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10240_ _03037_ _03119_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_131_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07528__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10200__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08944__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10171_ _02980_ _02988_ _03051_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_113_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06955__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13930_ _00261_ net101 clknet_leaf_19_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_89_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11700__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13861_ _00192_ net36 clknet_leaf_44_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_69_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12812_ _05577_ _05578_ _05588_ _05698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13792_ _00123_ net36 clknet_leaf_66_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_85_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10267__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12743_ _05530_ _05532_ _05624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07132__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12674_ _05508_ _05523_ _05548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_155_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11625_ _00378_ _01249_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11556_ _00387_ _01610_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07435__A2 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10507_ _03382_ _03383_ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11487_ _00384_ _01610_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11519__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13226_ _06056_ _06062_ _06147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10438_ _03221_ _03236_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07199__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13748__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13157_ _00375_ _03558_ _06072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10369_ _03239_ _03247_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06946__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10742__A2 _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12108_ _04950_ _04874_ _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13456__B _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13088_ _05994_ _05996_ _05997_ _05998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_53_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12039_ _00397_ _01693_ _04882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09360__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13920__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07580_ _00564_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10258__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09250_ _02060_ _02061_ _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08201_ net142 _05833_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09181_ _02070_ _02072_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ _01025_ _01033_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10430__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08063_ _00964_ _00963_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_71_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07014_ _05572_ _05452_ _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__09179__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13739__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06937__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11930__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08965_ _01834_ _01859_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07916_ _00803_ _00817_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08896_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[6\] _01792_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08154__A3 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07847_ _00737_ _00748_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13911__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07778_ DDS_Stage.xPoints_Generator1.RegFrequency\[-10\] DDS_Stage.xPoints_Generator1.RegF\[-10\]
+ _00402_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12238__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09517_ _02395_ _02405_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07114__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09448_ _02274_ _02336_ _02300_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08862__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09379_ _06664_ _00385_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09406__A3 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11410_ _04237_ _04250_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_124_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12390_ _05192_ _05201_ _05242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07417__A2 _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11341_ _04181_ _04182_ _04183_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_61_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11272_ _04111_ _04114_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08378__B1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13011_ _03189_ _00387_ _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10223_ _03095_ _03102_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_18_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11516__A4 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10154_ net61 net60 _06744_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_7_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10085_ _02965_ _02966_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10488__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13913_ _00244_ net36 clknet_leaf_53_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_89_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13902__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09893__A3 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13844_ _00175_ clknet_leaf_48_clk DDS_Stage.xPoints_Generator1.RegP\[-4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12229__A2 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13775_ _00110_ clknet_leaf_6_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07105__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10987_ _00372_ _02854_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12726_ _05517_ _05603_ _05604_ _05606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_85_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11452__A3 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12657_ _05362_ _05432_ _05531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11608_ _04446_ _04449_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07408__A2 _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12588_ _05369_ _05430_ _05454_ _05455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_41_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ _04381_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08081__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13209_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-6\] _06118_ _06128_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09030__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06919__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11912__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_146_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08750_ _00388_ _06618_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07701_ DDS_Stage.xPoints_Generator1.CosNew\[-1\] _00663_ _00577_ _00664_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08681_ _01577_ _01578_ _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07632_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-11\] _00604_ _00395_ _00605_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07563_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[5\] _00555_ _00395_ _00556_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_24_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09302_ _02111_ _02124_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07494_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-8\] _00499_ _00395_ _00500_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10246__A4 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10651__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ _02111_ _02124_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_146_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09164_ _02046_ _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10403__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08115_ _01003_ _01015_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09095_ _01985_ _01987_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10954__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ _00938_ _00939_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_61_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09021__A1 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDDS_Module_39 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_110_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07178__A4 _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09997_ _02869_ _02879_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08948_ _01757_ _01761_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09324__A2 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08879_ _01699_ _01701_ _01774_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_98_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10910_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-16\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-16\]
+ _05171_ _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07886__A2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11890_ _04700_ _04728_ _04730_ _04731_ _04732_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__07314__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10841_ _03704_ _03712_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07541__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13560_ _06457_ _06506_ _06507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_149_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _03643_ _03644_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08835__A1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12511_ _04012_ _04032_ _05371_ _05372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_109_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13491_ _06393_ _06432_ _06433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12442_ _04740_ _04741_ _05298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_87_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11198__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12373_ _05213_ _05219_ _05223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_22_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11324_ _04075_ _04093_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_127_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12147__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_29_clk_I clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11255_ _04096_ _04097_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09012__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10206_ _03086_ _03001_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11186_ _04026_ _04027_ _04028_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_128_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10137_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[21\] _03018_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13647__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09315__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10068_ _02948_ _02949_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07877__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12870__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10881__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13827_ _00158_ clknet_leaf_51_clk DDS_Stage.xPoints_Generator1.RegF\[-6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07451__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_48_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13758_ _00093_ clknet_leaf_58_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08826__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12709_ _05582_ _05586_ _05587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10633__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13689_ _00024_ clknet_leaf_2_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06862__I _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_61_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_44_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08054__A2 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09920_ _00373_ _06724_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09003__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12689__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09554__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09851_ _02718_ _02721_ _02735_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__11897__B1 _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08802_ _01612_ _01696_ _01697_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09782_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-11\] _02667_ _02668_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06994_ _06059_ _06632_ _06634_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08733_ _01628_ _01629_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_53_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11113__A2 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08664_ _01468_ _01469_ _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07615_ _00579_ _00588_ _00589_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08595_ _01489_ _01493_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_138_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ _05409_ _00541_ _06682_ _06146_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_37_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08817__A1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10624__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07477_ _05409_ _05995_ _06221_ _06787_ _06146_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09216_ _02106_ _02107_ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_146_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ _02024_ _02026_ _02039_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_17_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11719__A4 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09078_ _01770_ _01773_ _01863_ _01866_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__08596__A3 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ _05398_ _00385_ _00382_ _05833_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13867__CLK clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11040_ _03830_ _03831_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09545__A2 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07556__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11352__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13629__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10560__B1 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12991_ _05889_ _05890_ _05891_ _05892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_11942_ _04107_ _04784_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_123_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11873_ _04679_ _04688_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_129_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13612_ _06524_ _06561_ _06562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10824_ _03082_ _03695_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10615__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13543_ _06484_ _06487_ _06488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10755_ _03082_ _03600_ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__I1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13474_ _03556_ _00390_ _06414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10686_ _03401_ _03532_ _03559_ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12425_ _04105_ _05278_ _05279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_140_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12356_ _05194_ _05199_ _05205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_51_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11307_ net86 _02940_ _02938_ net83 _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12287_ _05068_ _05119_ _05129_ _05130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_11238_ _04078_ _04079_ _04080_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09536__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07446__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11343__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11169_ _03983_ _04011_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07462__B _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10854__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07400_ _00419_ _00420_ _00422_ _05182_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_63_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08380_ _00894_ _01279_ _01280_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07331_ _00375_ _00376_ _05182_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09472__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07262_ _05409_ _05691_ _05767_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09001_ _01838_ _01841_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07193_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-17\] _06804_ _05182_ _06805_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09224__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09224__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11031__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09903_ _02775_ _02786_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09527__A2 _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11334__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09834_ _02615_ _02618_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09765_ _00370_ _06710_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06977_ _06059_ _06617_ _06619_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13087__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ _01612_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11098__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09696_ _05182_ _02582_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer30 _05133_ net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
Xrebuffer41 net139 net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xrebuffer52 _02597_ net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_08647_ _01543_ _01544_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12047__B1 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08578_ _01399_ _01475_ _01476_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07529_ _05496_ _06806_ _05908_ _05658_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_76_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10073__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10540_ _05280_ net147 _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08018__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09215__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10471_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-3\] _03337_ _03347_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-2\]
+ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13011__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12210_ _05052_ _04946_ _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_121_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13190_ _06043_ _06107_ _06108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12141_ _04979_ _04983_ _04984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_124_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12117__A4 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12072_ _04893_ _04901_ _04915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07529__A1 _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11023_ _03863_ _03864_ _03865_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_60_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13078__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07282__B _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12974_ _05870_ _05871_ _05872_ _05873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_99_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10836__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11925_ _00365_ net135 _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11856_ _04675_ _04697_ _04698_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10807_ _05280_ _03679_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08257__A2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11787_ net54 _01693_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09454__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07304__I1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09454__B2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10738_ _03610_ _03538_ _03611_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13526_ _06467_ _06468_ _06470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_125_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13457_ _06322_ _06323_ _06325_ _06396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10669_ _00537_ _03540_ _03543_ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12408_ _05258_ _05260_ _05261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11013__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11013__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13388_ _00372_ _00375_ _03727_ _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12339_ _05154_ _05155_ _05145_ _05186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06900_ _05420_ _05463_ _05875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07880_ _00779_ _00780_ _00781_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__11867__A3 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09550_ _02360_ _02361_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_39_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12816__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08501_ net154 _01290_ _01400_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_76_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09481_ _02368_ _02369_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08496__A2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11095__A4 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08432_ _01331_ _01237_ _01233_ _01235_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ _06308_ _00388_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08248__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09445__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13241__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07314_ _00361_ net60 _05182_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08294_ _01173_ _01192_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_34_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07245_ _05518_ _06211_ _06732_ _05409_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_27_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07176_ _06726_ _06789_ _06790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11555__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08420__A2 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11307__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09817_ net95 _06679_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09920__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07931__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07931__B2 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09748_ _02555_ _02556_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09679_ _02453_ _02454_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11710_ _04549_ _04551_ _04552_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12690_ net86 net84 _03679_ _03725_ _05566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_84_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08418__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11641_ _04482_ _04483_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_154_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12035__A3 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09987__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11572_ _00384_ _01247_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13311_ _05953_ _05959_ _06152_ _06238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__07998__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10523_ _03138_ _03309_ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput19 net100 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_134_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13242_ _00372_ _03725_ _06164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06960__I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ _03249_ _03252_ _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_122_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13173_ _03266_ _00390_ _06089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10385_ _03257_ _03262_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_131_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12124_ _00361_ _02499_ _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13299__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12055_ _04895_ _04896_ _04898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08175__A1 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11006_ _03792_ _03794_ _03848_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07922__A1 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__B1 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12957_ _05801_ _05816_ _05855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11908_ _04749_ _04750_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12888_ _05682_ _05779_ _05780_ _05781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11839_ net66 net54 _01524_ _01430_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_28_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10037__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07989__A1 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07989__B2 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13509_ _06439_ _06449_ _06450_ _06451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_125_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07030_ _05822_ _06664_ _06665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11537__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08981_ _01805_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_71_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07932_ _00832_ _00833_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_71_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07863_ _06618_ _00370_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09602_ _02487_ _02393_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07794_ DDS_Stage.xPoints_Generator1.RegFrequency\[-2\] DDS_Stage.xPoints_Generator1.RegF\[-2\]
+ _00402_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09533_ _02356_ _02364_ _02420_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_149_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11473__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10276__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09464_ net137 _06730_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07141__A2 _06759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08415_ _00981_ _01244_ _01315_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09395_ _02280_ _02284_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_47_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08346_ _05280_ _01247_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12973__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08277_ _01177_ _01178_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07228_ _05387_ _00292_ _00293_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07159_ _05387_ _06773_ _06775_ _06776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_113_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10200__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _02983_ _03050_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08157__A1 _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11700__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13860_ _00191_ net36 clknet_leaf_48_clk DDS_Stage.xPoints_Generator1.RegFrequency\[-3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_12811_ _05696_ _05587_ _05697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_2_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13791_ _00122_ net36 clknet_leaf_73_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_97_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10267__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12742_ _05619_ _05622_ _05623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_69_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12673_ _05508_ _05523_ _05547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_139_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11624_ _00372_ _00375_ _01524_ _01430_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_65_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11216__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06891__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11555_ _00381_ _01792_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10506_ _03209_ _03289_ _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11486_ _04217_ _04327_ _04328_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11519__A2 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13225_ _06079_ _06102_ _06144_ _06145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10437_ _03274_ _03314_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13156_ _03556_ _00378_ _06071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10368_ _03082_ _03246_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__06946__A2 _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12107_ _00381_ _00384_ _02051_ _01956_ _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_13087_ net147 _00381_ _05997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10299_ _03175_ _03176_ _03177_ _03178_ _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__08148__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12038_ _04877_ _04880_ _04881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09896__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_144_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09648__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_29_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11455__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10258__A2 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08200_ net60 net73 _05833_ _05398_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_146_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06882__A1 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09180_ _01999_ _02000_ _02071_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08131_ _01028_ _01032_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09820__A1 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08062_ _00774_ _00783_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10430__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12707__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07013_ _06059_ _06648_ _06650_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08387__A1 _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06937__A2 _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11930__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08964_ _01842_ _01858_ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08139__A1 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07915_ _00811_ _00816_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08895_ _01784_ _01790_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11143__B1 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone6_I net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07846_ _00742_ _00747_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08154__A4 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09639__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ _00704_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09516_ _01967_ _02398_ _02404_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_84_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09447_ _02202_ _02218_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08862__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06873__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09378_ _06659_ _00388_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12946__A1 _05740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08329_ _01173_ _01192_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09406__A4 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11340_ _00387_ _01249_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11271_ _04039_ _04113_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13010_ _05810_ _05911_ _05912_ _05913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08378__A1 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08378__B2 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10222_ _03095_ _03102_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_30_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10185__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07050__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _02608_ _02704_ _03033_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_7_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10084_ _00398_ _00394_ _06685_ _06691_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__07274__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09878__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13912_ _00243_ net36 clknet_leaf_54_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__10488__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11685__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08550__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09893__A4 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13843_ _00174_ clknet_leaf_49_clk DDS_Stage.xPoints_Generator1.RegP\[-5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10986_ _03828_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13774_ _00109_ clknet_leaf_15_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08302__A1 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12725_ _05519_ _05520_ _05604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_29_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11452__A4 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06864__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12656_ _05528_ _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11607_ _04446_ _04449_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12587_ _05372_ _05429_ _05454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11538_ _00378_ _01794_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11469_ _00361_ _00365_ _02153_ _02051_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_111_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13208_ _06029_ _06121_ _06127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09030__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10176__A1 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11912__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13139_ _05978_ _06001_ _06051_ _06052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_146_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07592__A2 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13114__A1 _06021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07700_ DDS_Stage.xPoints_Generator1.RegFrequency\[-1\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-1\]
+ _00662_ _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_40_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08680_ _06308_ _00398_ _00394_ net153 _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_07631_ DDS_Stage.xPoints_Generator1.CosNew\[-11\] _00603_ _00577_ _00604_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07562_ _05409_ _00541_ _06693_ _05658_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_24_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09301_ _02174_ _02177_ _02191_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_66_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07493_ _06790_ _06827_ _00455_ _06797_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09232_ _02115_ _02123_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_150_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09163_ _01513_ _01518_ _02054_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_56_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08114_ _01003_ _01015_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11600__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09094_ _01898_ _01899_ _01986_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ _00946_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_141_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09021__A2 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07032__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09996_ _02876_ _02878_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_86_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08947_ _01835_ _01838_ _01841_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_99_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08878_ _01770_ _01773_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__13896__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07829_ _06308_ _00379_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07886__A3 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10840_ _03706_ _03711_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11419__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10771_ _00394_ _06744_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08835__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06846__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12510_ _03982_ _05370_ _04011_ _05371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13490_ _06407_ _06431_ _06432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12441_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-23\] _05296_ _05297_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08599__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11198__A3 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12372_ _05211_ _05221_ _05222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_97_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11323_ _04094_ _04162_ _04163_ _04164_ _04165_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__07271__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13344__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12147__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11254_ _03853_ _03913_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13287__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09012__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10205_ _02945_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11185_ _02854_ _00381_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08771__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ _03017_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_128_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13647__A2 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10067_ _02880_ _02888_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09315__A3 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13887__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10330__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12870__A3 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13826_ _00157_ clknet_leaf_51_clk DDS_Stage.xPoints_Generator1.RegF\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13757_ _00092_ clknet_leaf_59_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08826__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _03795_ _03798_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_127_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12708_ _05584_ _05585_ _05586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10633__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13688_ _00023_ clknet_leaf_2_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12639_ _02762_ _00390_ _05511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_139_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_139_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08054__A3 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09251__A2 _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13811__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07262__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13335__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09003__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07014__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ _02726_ _02734_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08801_ _01616_ _01686_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06993_ _05822_ _06633_ _06634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09781_ _02501_ _02574_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08732_ _06654_ _00370_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13878__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08663_ _01468_ _01469_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10321__A1 _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07614_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-14\] DDS_Stage.xPoints_Generator1.RegFrequency\[-14\]
+ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08594_ _01490_ _01491_ _01492_ _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_49_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12074__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13660__B _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07545_ _05572_ _05550_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08817__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10624__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07476_ _05658_ _00484_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09215_ _06637_ _00394_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ _02030_ _02038_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_60_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10388__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13802__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07253__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09077_ _01776_ _01778_ _01779_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08596__A4 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13326__A1 _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ _00929_ _00768_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_13_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07005__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07800__I0 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10560__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09979_ _02822_ _02831_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13629__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10560__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12990_ _03556_ _00372_ _05891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13869__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11941_ _04783_ _04108_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10312__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11872_ _04712_ _04714_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13611_ _06553_ _06560_ _06561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_156_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10823_ _03401_ _03694_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13542_ _06485_ _06486_ _06487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10754_ _03551_ _03622_ _03624_ _03625_ _03626_ _03545_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_0_82_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10685_ _03082_ _03533_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13473_ _03485_ _00393_ _06413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12424_ _04174_ _05276_ _05277_ _05278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07244__A1 _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12355_ _05192_ _05201_ _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06912__B _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13317__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11306_ _00359_ _02854_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12286_ _05121_ _05122_ _05128_ _05129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_50_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11237_ net87 net83 _03018_ _02940_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_11168_ _03999_ _04010_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10551__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10119_ _02992_ _03000_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11099_ net84 _03416_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10303__A1 _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10854__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13809_ _00140_ net36 clknet_leaf_66_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_63_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_60_clk_I clknet_3_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07330_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-8\] _00376_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11803__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09472__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07483__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ _00320_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09000_ _01838_ _01841_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_75_clk_I clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07192_ _05658_ _06802_ _06803_ _06715_ _06804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__09224__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07235__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11031__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08983__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09902_ _02783_ _02785_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09833_ _02632_ _02640_ _02717_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_13_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09764_ _02647_ _02649_ _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06976_ _05822_ _06618_ _06619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08715_ _01602_ _01604_ _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11098__A2 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09695_ _02575_ _02580_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer20 _00964_ net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer42 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-15\] net141 vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10845__A2 _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08646_ _06637_ _00373_ _01462_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_68_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12047__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_28_clk_I clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12047__B2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08577_ _01401_ _01415_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07528_ _05409_ _06715_ _06566_ _06146_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_92_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__A2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07459_ _05658_ _00469_ _00470_ _06711_ _05182_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__07474__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13547__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10470_ _03328_ _03335_ _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_33_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09215__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07226__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09129_ _02020_ _02021_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12140_ _04982_ _04983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10781__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12071_ _04887_ _04905_ _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11022_ _03858_ _03862_ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12973_ _00361_ _03725_ _05872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11924_ _00361_ _02586_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11855_ _04645_ _04674_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_72_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold92_I Enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10806_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[29\] _03679_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_45_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11786_ net66 _01792_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09454__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10429__B _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13525_ _06463_ _06464_ _06466_ _06468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_55_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07465__A1 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10737_ _03539_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13456_ _06239_ _06328_ _06237_ _06395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10668_ _03541_ _03542_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12407_ _05259_ _04172_ _05260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11013__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13387_ _06249_ _06250_ _06248_ _06321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10599_ _03333_ _03473_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12338_ _05178_ _05183_ _05184_ _05185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_10_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_81_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12269_ _05093_ _05098_ _05111_ _05112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11867__A4 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09142__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08500_ _01281_ _01285_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09480_ _02200_ _02298_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_90_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08431_ _00983_ _01329_ _01330_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08362_ _06523_ _00382_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09445__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07313_ _00362_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_16
XANTENNA__07456__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08293_ _01070_ _01071_ _01073_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_46_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13529__A1 _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07244_ _00305_ _00306_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07208__B2 _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07175_ _05420_ _05485_ _05409_ _06789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_76_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09816_ _02696_ _02700_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07931__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_129_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09747_ _02555_ _02556_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_20_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06959_ _06146_ _06502_ _06513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09678_ _00373_ _06696_ _02455_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_120_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08629_ _01509_ _01433_ _01507_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_96_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11640_ _04416_ _04419_ _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12035__A4 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11571_ _00381_ _01249_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13310_ _05953_ _06152_ _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__07998__A2 _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10522_ _03295_ _03397_ _03398_ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_134_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_138_Left_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_118_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13241_ _00375_ _03679_ _06163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10453_ _03249_ _03252_ _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13172_ _03189_ _00393_ _06088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10384_ _03257_ _03262_ _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12123_ _00369_ _02238_ _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12054_ _04895_ _04896_ _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08175__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11005_ _03815_ _03846_ _03847_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07922__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__B2 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12956_ _05751_ _05819_ _05853_ _05854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_99_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11907_ _00381_ _02236_ _02153_ _00384_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_87_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12887_ _05683_ _05684_ _05780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_114_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11838_ net66 _01524_ _01430_ net54 _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_114_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10159__B _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07438__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11769_ _04609_ _04610_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_138_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07989__A2 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13508_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-2\] _06446_ _06448_ _06450_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_82_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13439_ _06363_ _06376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_58_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07610__A1 _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ _01795_ _01874_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07931_ _05864_ _00388_ _00385_ _06179_ _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_71_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07862_ _00736_ _00763_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09601_ _02055_ _02062_ _02488_ _02138_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_07793_ _00712_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09115__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09532_ _02342_ _02355_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09463_ net96 _06659_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11473__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08414_ _00930_ _00980_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09394_ _02281_ _02282_ _02283_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_19_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07429__A1 _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08345_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[0\] _01247_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__12422__A1 _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_clk clknet_3_5__leaf_clk clknet_leaf_31_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12973__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ _01175_ _01176_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ _05182_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-11\] _00293_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ _06092_ _06774_ _06757_ _06146_ _06775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_113_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07089_ _06713_ _06714_ _06715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_113_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12489__A1 _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08157__A2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11161__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11700__A3 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12810_ _05581_ _05696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_2_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13790_ _00121_ net36 clknet_leaf_62_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_2_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12741_ _05453_ _05620_ _05621_ _05622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12672_ _05461_ _05526_ _05545_ _05546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_146_Left_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11623_ _04464_ _04465_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06891__A2 _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11216__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_22_clk clknet_3_6__leaf_clk clknet_leaf_22_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_41_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08093__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11554_ _00384_ _01693_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10975__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10505_ _03285_ _03288_ _03382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07288__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11485_ _04215_ _04216_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13224_ _06055_ _06078_ _06144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold55_I FreqPhase[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10436_ _03292_ _03313_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10727__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13155_ _05955_ _06067_ _06068_ _06069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10367_ _03242_ _03245_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12106_ _04948_ _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_155_Left_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13086_ _03340_ _00384_ _05996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10298_ _02842_ _02843_ _02844_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__08148__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12037_ _04743_ _04879_ _04880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11152__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09896__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09648__A2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11455__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12939_ _05629_ _05831_ _05837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13_clk clknet_3_6__leaf_clk clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08130_ _01029_ _01030_ _01031_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_16_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10966__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08061_ _00953_ _00961_ _00962_ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10430__A3 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07012_ _05822_ _06649_ _06650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12707__A2 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10718__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08387__A2 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09584__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11930__A3 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08963_ _01844_ _01857_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08139__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07914_ _00812_ _00815_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08894_ _01787_ _01789_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11143__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11143__B2 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07845_ _00743_ _00746_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13663__B _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclone5 _02607_ net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07776_ DDS_Stage.xPoints_Generator1.RegFrequency\[-11\] DDS_Stage.xPoints_Generator1.RegF\[-11\]
+ _00402_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09639__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09515_ _02399_ _02403_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09446_ _02333_ _02334_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06873__A2 _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09377_ _00382_ _06672_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08328_ _01215_ _01225_ _01228_ _01229_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_117_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07822__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ _01155_ _01160_ _05398_ _00370_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_115_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11270_ _04112_ _04040_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08378__A2 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10221_ _02931_ _03096_ _03098_ _03099_ _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__10185__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10152_ net63 _06701_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07050__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10083_ _00398_ _06685_ _06691_ _00394_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09878__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13911_ _00242_ net36 clknet_leaf_53_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07889__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11685__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08550__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13842_ _00173_ clknet_leaf_49_clk DDS_Stage.xPoints_Generator1.RegP\[-6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13773_ _00108_ clknet_leaf_15_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10985_ _00378_ _02586_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08302__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12724_ _05519_ _05520_ _05603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06864__A2 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12655_ _05453_ _05455_ _05527_ _05528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_53_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11606_ _04447_ _04448_ _04226_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_12586_ _05451_ _05368_ _05453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10948__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11537_ _00372_ _02051_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11468_ _00361_ _02153_ _02051_ _00365_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_150_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13207_ _05822_ _06124_ _06126_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09566__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10419_ _03126_ _03211_ _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11373__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11399_ net87 _02238_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10176__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13138_ _05952_ _05977_ _06051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_146_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09318__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13069_ _05961_ _05976_ _05977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_clk clknet_3_2__leaf_clk clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12873__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07630_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-11\] DDS_Stage.xPoints_Generator1.RegFrequency\[-11\]
+ _00602_ _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_88_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12625__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07561_ _06059_ _00552_ _00553_ _00554_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_49_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09300_ _02182_ _02190_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_24_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07492_ _00495_ _00497_ _00498_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07701__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09231_ _02118_ _02122_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_146_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08057__A1 _06523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09162_ _01700_ _02053_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__13050__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08113_ _01006_ _01014_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_114_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11600__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09093_ _06664_ _00373_ _01900_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_32_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ _00942_ _00943_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07280__A2 _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09021__A3 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09995_ _02608_ _02704_ _02877_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__09309__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08946_ _01839_ _01840_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08877_ _01619_ _01771_ _01772_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07828_ net155 _00373_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07886__A4 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11419__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07759_ _00695_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10627__B1 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10770_ _00398_ _06742_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07343__I0 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09429_ _02306_ _02309_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08048__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12440_ _05190_ _05295_ _05296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08599__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12371_ _05213_ _05219_ _05220_ _05221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__11198__A4 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11322_ _04076_ _04089_ _04162_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_132_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13344__A2 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11253_ _04075_ _04093_ _04095_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10204_ _03022_ _03025_ _03084_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_11184_ _02762_ _00384_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08771__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10135_ _02940_ _03016_ _00395_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_128_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10066_ _02869_ _02879_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09315__A4 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09720__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10330__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12870__A4 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13825_ _00156_ clknet_leaf_51_clk DDS_Stage.xPoints_Generator1.RegF\[-8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12607__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13756_ _00091_ clknet_leaf_59_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10968_ _03807_ _03810_ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_106_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10094__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12707_ _03340_ _00372_ _05585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13687_ _00022_ clknet_leaf_0_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10899_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-21\] _03765_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12638_ _02586_ _00393_ _05510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12569_ _03971_ _04035_ _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08054__A4 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09539__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13335__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07014__A2 _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08800_ _01616_ _01686_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09780_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-10\] _02659_ _02665_ _02666_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06992_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-15\] _06633_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08731_ _01624_ _01627_ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08662_ _01556_ _01559_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07613_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-14\] DDS_Stage.xPoints_Generator1.RegFrequency\[-14\]
+ _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08593_ net60 _06654_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07544_ _05387_ _00537_ _00538_ _00540_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__12074__A2 _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07475_ _06651_ _06373_ _06754_ _06756_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clone22_I net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09214_ _06633_ _00398_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09145_ _02033_ _02037_ _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_101_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11585__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10388__A2 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13388__B _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09076_ _01968_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_79_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07253__A2 _06623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08027_ _00928_ _00869_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_102_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08202__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09950__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09978_ _02772_ _02821_ _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10560__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08929_ _01731_ _01732_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_110_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11940_ _00381_ _00384_ _02238_ _02236_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_54_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11871_ _00361_ _01247_ _04713_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_54_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13610_ _06556_ _06559_ _06560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_10822_ _03693_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08269__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13541_ _00390_ _03558_ _06486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10753_ _03544_ _03546_ _03616_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_82_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13472_ net147 _00397_ _06412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10684_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[28\] _03558_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_125_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12423_ _04106_ _04173_ _05277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_51_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12354_ _05192_ _05201_ _05202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_106_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13317__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06912__C _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11305_ _04128_ _04129_ _04130_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07296__B _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12285_ _05124_ _05127_ _05128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11236_ net87 _03018_ _02940_ net84 _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10000__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11167_ _04000_ _04009_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10118_ _02998_ _02999_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11098_ _00351_ _03485_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10049_ _02758_ _02850_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07180__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13808_ _00139_ net36 clknet_leaf_66_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_19_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13739_ _00074_ net36 clknet_leaf_73_clk DDS_Stage.xPoints_Generator1.CosNew\[-14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__11803__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13005__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07260_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-5\] _00319_ _00320_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_14_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08680__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__A2 _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07191_ _05658_ _06681_ _06803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07235__A2 _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13796__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08983__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06994__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12516__B1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09901_ _02608_ _02704_ _02784_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09832_ _02635_ _02639_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10542__A2 _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09763_ _02547_ _02548_ _02648_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06975_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-17\] _06618_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08714_ _06059_ _01609_ _01611_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09694_ _02575_ _02580_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xrebuffer10 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-14\] net62 vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xrebuffer21 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-13\] net90 vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
Xrebuffer32 _00391_ net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08645_ _01460_ _01461_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07171__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12047__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08576_ _01401_ _01415_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09999__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07527_ _05387_ _00522_ _00526_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07458_ _05658_ _00451_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13547__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07389_ DDS_Stage.xPoints_Generator1.CosNew\[-3\] DDS_Stage.xPoints_Generator1.RegP\[-3\]
+ _00402_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _06633_ _00394_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07226__A2 _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13787__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ _01798_ _01867_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_124_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12070_ _04907_ _04910_ _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_124_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11021_ _03822_ _03823_ _03825_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_60_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12972_ _00365_ _03679_ _05871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13483__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11923_ _00369_ _02499_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07162__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11854_ _04694_ _04695_ _04696_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__10049__A1 _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10805_ _05182_ _03677_ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11785_ _04625_ _04626_ _04627_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13524_ _06463_ _06464_ _06466_ _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_hold85_I FreqPhase[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10736_ _03541_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_137_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13455_ _06331_ _06355_ _06392_ _06393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10667_ _03476_ _03479_ _03472_ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12406_ _04141_ _04145_ _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13386_ _06239_ _06253_ _06237_ _06320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10598_ _03473_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12337_ _05180_ _05181_ _05184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06976__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12268_ _05096_ _05097_ _05111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11219_ _04059_ _04060_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12199_ _00372_ _00375_ _02153_ _02051_ _05042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13950__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13474__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09142__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07153__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08430_ _01069_ _01094_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06900__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08361_ _00913_ _01260_ _01261_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08102__B1 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07312_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-12\] _00362_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08292_ _01171_ _01193_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07456__A2 _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-8\] _00306_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07174_ _05409_ _05875_ _06788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09905__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11712__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09815_ _02697_ _02698_ _02699_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__13941__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09746_ _02628_ _02631_ _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06958_ _06447_ _06469_ _06491_ _06502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09677_ _02448_ _02466_ _02563_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06889_ _05658_ _05724_ _05745_ _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_68_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ _01510_ _01519_ _01508_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_87_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13217__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08559_ _01371_ _01456_ _01457_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11570_ _04224_ _04412_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_76_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07447__A2 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10521_ _03298_ _03312_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07998__A3 _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13240_ _00378_ _03558_ _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10452_ _03329_ _03253_ _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13171_ _03018_ _00397_ _06087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10383_ _03102_ _03258_ _03261_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12122_ _04960_ _04964_ _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12053_ _00365_ _02499_ _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11703__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11004_ _03835_ _03845_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13932__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13456__A1 _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_74_clk_I clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__A2 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12955_ _05753_ _05818_ _05853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07135__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11906_ _00381_ _00384_ _02236_ _02153_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_12886_ _05683_ _05684_ _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11837_ net70 _01249_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11768_ _04609_ _04610_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_126_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10719_ _03589_ _03592_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13507_ _06446_ _06448_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-2\] _06449_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11699_ net66 _01792_ _01693_ net54 _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_24_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_clk_I clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13438_ _06304_ _06361_ _06375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xrebuffer1 _02754_ net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10890__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13369_ _06204_ _06208_ _06290_ _06301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_51_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06949__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_27_clk_I clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07930_ _06179_ _05864_ _00388_ _00385_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_139_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07861_ _00749_ _00762_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13923__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09600_ _02227_ _02487_ _02393_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_07792_ DDS_Stage.xPoints_Generator1.RegFrequency\[-3\] DDS_Stage.xPoints_Generator1.RegF\[-3\]
+ _00402_ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09115__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09531_ _02340_ _02417_ _02418_ _02365_ _02386_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__07126__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09462_ _00355_ _06724_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08413_ _01310_ _01313_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09393_ net142 _06701_ _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08344_ _00981_ _01244_ _05182_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08626__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07429__A2 _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08275_ _01175_ _01176_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_73_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer32_I _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07226_ _05658_ _06681_ _06830_ _06831_ _06796_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_116_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12186__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07157_ _05409_ _06726_ _06774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07088_ _05420_ _06070_ _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_113_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13914__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11161__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11700__A4 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A2 _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _02525_ _02613_ _02614_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_2_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07117__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12740_ _05455_ _05527_ _05621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12671_ _05465_ _05525_ _05545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_93_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11622_ _04289_ _04342_ _04225_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__10424__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11553_ _04332_ _04394_ _04395_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08093__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10975__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10504_ _03306_ _03311_ _03380_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_133_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11484_ _04215_ _04216_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13223_ _06141_ _06142_ _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10435_ _03295_ _03298_ _03312_ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_27_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11924__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13154_ _05956_ _05957_ _06068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_0_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10366_ _03243_ _03244_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12105_ _04945_ _04946_ _04947_ _04948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13085_ _03266_ _00387_ _05994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10297_ _02839_ _02493_ _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_109_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12036_ _04878_ _04744_ _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_53_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13905__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11152__A2 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07108__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09648__A3 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08856__A1 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12938_ _05720_ _05722_ _05836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12869_ net54 _03725_ _03727_ net66 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07479__B _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09820__A3 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10966__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08060_ _00957_ net85 _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07011_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-12\] _06649_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_141_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09584__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08962_ _01848_ _01856_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11930__A4 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07913_ _00813_ _00814_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08893_ _01788_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11143__A2 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07844_ _00744_ _00745_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07775_ _00703_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclone6 net59 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_151_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09514_ _02314_ _02401_ _02402_ _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_78_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09445_ _00370_ _06696_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09376_ _02186_ _02264_ _02265_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10406__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08327_ _01219_ _01223_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_145_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08258_ _01147_ _01157_ _01158_ _01159_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07822__A2 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07209_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-14\] _06817_ _05182_ _06818_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09024__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08189_ _01085_ _01090_ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11906__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10220_ _02673_ _02675_ _02680_ _03100_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_104_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10151_ _02954_ _02959_ _03031_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13659__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10082_ _02704_ _02962_ _02963_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13910_ _00241_ net36 clknet_leaf_54_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07889__A2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13841_ _00172_ clknet_leaf_51_clk DDS_Stage.xPoints_Generator1.RegP\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13772_ _00107_ clknet_leaf_10_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10984_ _03824_ _03825_ _03826_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10645__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12723_ _05598_ _05601_ _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_128_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12654_ _05461_ _05526_ _05527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11605_ net86 _02153_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09263__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12585_ _05365_ _05451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10948__A2 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11536_ _00375_ _01956_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07274__B1 _06759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11467_ _04280_ _04308_ _04309_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_80_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13206_ _05280_ net34 _06126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10418_ _03207_ _03210_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09566__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11398_ net84 _02236_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11373__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__B1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13137_ _06046_ _06049_ _06050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10349_ _03147_ _03148_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09318__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13068_ _05965_ _05975_ _05976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12019_ _04855_ _04856_ _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12873__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07560_ _05409_ _05594_ _06735_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12625__A2 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07491_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-9\] _00498_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09230_ _02119_ _02120_ _02121_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_119_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09161_ _01774_ _01867_ _01947_ _02047_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_57_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13050__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08112_ _01009_ _01013_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_71_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11061__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09092_ _01893_ _01983_ _01984_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_4_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08043_ _00942_ _00943_ _00944_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_71_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09021__A4 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ net63 _06691_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09309__A2 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08945_ _00398_ _00394_ _06598_ _06618_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_08876_ _01622_ _01684_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10875__A1 _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07827_ _06059_ _00575_ _00729_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07758_ net110 DDS_Stage.xPoints_Generator1.RegP\[-5\] _00684_ _00695_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10627__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10627__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ _00653_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07343__I1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _02317_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10538__B _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09359_ _02246_ _02248_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__08048__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12370_ _05217_ _05218_ _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_63_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11321_ _04121_ _04139_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_90_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07339__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11252_ _04090_ _04094_ _04092_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10203_ _03072_ _03083_ _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11183_ _00387_ _02586_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10134_ _03013_ _03015_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_128_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10065_ _02890_ _02911_ _02946_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09720__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10330__A3 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13824_ _00155_ clknet_leaf_68_clk DDS_Stage.xPoints_Generator1.RegF\[-9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12607__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11815__B1 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13755_ _00090_ clknet_leaf_59_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10967_ _03808_ _03809_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09484__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12706_ _03266_ _00375_ _05584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10094__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10898_ _05387_ _03763_ _03764_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13686_ _00021_ clknet_leaf_1_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07601__I _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12637_ net135 _00397_ _05509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_139_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12568_ _03977_ _05433_ _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_136_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_152_Right_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11519_ _00351_ _02584_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12499_ _05356_ _05359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07249__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09539__A2 _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06991_ _05658_ _06631_ _06632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08730_ _01625_ _01626_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08661_ _01557_ _01558_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07612_ _00584_ _00587_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08592_ net91 _06649_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07712__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07543_ _05182_ _00539_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07474_ _06059_ _00482_ _00483_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09213_ _02027_ _02103_ _02104_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09227__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09144_ _02034_ _02035_ _02036_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12782__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11585__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09075_ _01943_ _01946_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_79_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08450__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08026_ _00927_ _00876_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_130_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08202__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09977_ _02858_ _02859_ _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08928_ _01731_ _01732_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_118_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08859_ net60 _06664_ _06659_ net61 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11870_ _04707_ _04711_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_123_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10821_ _03691_ _03692_ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08269__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13540_ _03556_ _00393_ _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11273__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10752_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[2\] _03623_ _03625_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_149_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13471_ _06244_ _06326_ _06410_ _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10683_ _03553_ _03555_ _03557_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12422_ _05250_ _05270_ _05275_ _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11025__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12353_ _05194_ net82 _05200_ _05201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_2_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11304_ _04127_ _04135_ _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12284_ _04954_ _05125_ _05126_ _05127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12525__A1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11235_ _00359_ _02938_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11166_ _04003_ _04008_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07952__A1 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _00370_ _06742_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11097_ _00359_ _03340_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10048_ _02849_ _02930_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07704__A1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold90 LoadP net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_117_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13807_ _00138_ net36 clknet_leaf_66_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_129_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09457__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11999_ _04840_ _04841_ _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_63_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11264__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13738_ _00073_ net36 clknet_leaf_73_clk DDS_Stage.xPoints_Generator1.CosNew\[-15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_128_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11803__A3 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13005__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13669_ _00004_ clknet_leaf_78_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08680__A2 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__A3 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11016__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07190_ _05409_ _05550_ _05691_ _06802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_131_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07487__B _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07235__A3 _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12516__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09900_ net95 _06685_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12516__B2 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08196__A1 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09831_ _02691_ _02707_ _02715_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__07943__A1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06974_ _05658_ _06616_ _06617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09762_ _00373_ _06701_ _02549_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08713_ _05280_ _01610_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09693_ _02576_ _02577_ _02579_ _02405_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09696__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer11 _00960_ net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xrebuffer22 _00366_ net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08644_ _01455_ _01473_ _01541_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xrebuffer33 net96 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_83_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xrebuffer55 _01286_ net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_89_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08575_ _01455_ _01473_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_117_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer62_I net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07526_ _05658_ _00524_ _00525_ _00330_ _05171_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__09999__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08120__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07457_ _05431_ _06705_ _00468_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_134_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07388_ _00414_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09127_ _00398_ _06627_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09058_ _00449_ _01947_ _01951_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_102_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08009_ _00831_ _00832_ _00833_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_130_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13180__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07617__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11020_ _03858_ _03862_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_124_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12971_ _00369_ _03558_ _05870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13483__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11494__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11922_ _04760_ _04764_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12691__B1 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11853_ _04651_ _04670_ _04671_ _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_10804_ _03627_ _03675_ _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_103_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11784_ net66 net54 _01693_ _01610_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_103_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13523_ _06409_ _06430_ _06465_ _06466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_31_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10735_ _03605_ _03608_ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_125_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10666_ _03468_ _03471_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13454_ _06320_ _06329_ _06392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07870__B1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12405_ _04866_ _05251_ _05256_ _05257_ _05258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_13385_ _06256_ _06281_ _06317_ _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10597_ _03328_ _03410_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_152_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12336_ _05180_ _05181_ _05183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06976__A2 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12267_ _05051_ _05054_ _05109_ _05110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__13171__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11218_ _04059_ _04060_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_12198_ _00378_ _01956_ _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11149_ _03989_ _03990_ _03991_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__10888__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09678__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13474__A2 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07153__A2 _06765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06900__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08360_ _00914_ _00915_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_53_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11237__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08102__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07311_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-12\] _00361_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
XANTENNA__08102__B2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08291_ _01173_ _01192_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_46_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07242_ _00302_ _00303_ _00304_ _05182_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_144_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07173_ _05420_ _05886_ _06787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_76_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08169__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09905__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11712__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09814_ net60 _06738_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_107_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09745_ _02629_ _02630_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06957_ _06232_ _06480_ _06081_ _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_94_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09669__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06888_ _05409_ _05734_ _05745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09676_ _02451_ _02465_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_68_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_6_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08627_ _01522_ _01523_ _01525_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_87_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13217__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08558_ _01395_ _01398_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07509_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-5\] _00512_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08489_ _01369_ _01388_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_147_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10520_ _03298_ _03312_ _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_130_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07998__A4 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12728__A1 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10451_ _03170_ _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_118_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13170_ _06084_ _05972_ _06085_ _06086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11400__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10382_ _03259_ _03260_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12121_ _04961_ _04963_ _04964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07080__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07347__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12052_ _00361_ _02584_ _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07907__A1 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11703__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ _03835_ _03845_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07590__B _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12954_ _05748_ _05749_ _05747_ _05852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11905_ _00387_ _02051_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12885_ _05759_ _05776_ _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06894__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11836_ _04676_ _04678_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07810__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11767_ _04509_ _04510_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13506_ _06375_ _06377_ _06437_ _06448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_10718_ _03311_ _03591_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__07843__B1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11698_ net70 _01610_ _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12719__A1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13437_ _06298_ _06374_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10649_ _00382_ _03522_ _03523_ _03388_ _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_24_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer2 _04155_ net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13368_ _06291_ _06288_ _06299_ _06300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_58_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07071__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12319_ _05130_ _05163_ _05164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__07071__B2 _06698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13299_ _03189_ _00397_ _06182_ _06225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13144__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07860_ _00756_ _00760_ _00761_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07791_ _00711_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09530_ _02356_ _02364_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06895__I _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07126__A2 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09461_ _02345_ _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_149_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08412_ _00768_ _01311_ _01312_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__06885__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09392_ net92 _06696_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07720__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08343_ _00981_ _01244_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09823__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08626__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08274_ net152 _00370_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11630__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07225_ _06232_ _06211_ _06756_ _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_15_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer25_I _05740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12186__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07156_ _05658_ _06766_ _06772_ _06773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07062__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07087_ _05572_ _05550_ _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_112_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13135__A1 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07989_ _00363_ _06633_ _06627_ net91 _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09728_ _02526_ _02527_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07117__A2 _06737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09659_ _00373_ _06701_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06876__A1 _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12670_ _05458_ _05460_ _05544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_139_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11621_ _04440_ _04462_ _04463_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_38_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09814__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10424__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11552_ _00381_ _00384_ _01693_ _01610_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_37_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08093__A3 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10503_ _03301_ _03379_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13850__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10975__A3 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11483_ _04273_ _04282_ _04325_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_21_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10434_ _03306_ _03311_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_13222_ _06136_ _06137_ _06140_ _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_21_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11924__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07053__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13153_ _05956_ _05957_ _06067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10365_ _03138_ _03141_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13126__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12104_ _00381_ _00384_ _01956_ _01794_ _04947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_13084_ _05914_ _05991_ _05992_ _05993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10296_ _02839_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_97_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12035_ _00381_ _00384_ _02153_ _02051_ _04878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_53_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11688__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_144_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09648__A4 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12937_ _05443_ _05832_ _05835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_34_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08856__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06867__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12868_ _05668_ _05673_ _05758_ _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11819_ net54 _01610_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12799_ net147 _00372_ _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07010_ _06146_ _06647_ _06648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_70_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13365__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07044__A1 _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07595__A2 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08961_ _01851_ _01855_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07912_ _00391_ _05398_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11679__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08892_ _01529_ _01689_ _01688_ _01690_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_87_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07843_ _05833_ _00388_ _00385_ _05864_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07774_ DDS_Stage.xPoints_Generator1.RegFrequency\[-12\] DDS_Stage.xPoints_Generator1.RegF\[-12\]
+ _00402_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclone7 net88 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_79_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-14\] _02400_ _02402_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_78_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10103__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09444_ _02330_ _02332_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_66_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _02187_ _02188_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_148_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_96_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10406__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08326_ _01177_ _01226_ _01227_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_34_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08257_ net73 _05864_ _01148_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07283__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07208_ _06362_ _06768_ _06816_ _06761_ _06817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_115_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08188_ _01053_ _01089_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_73_clk_I clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09024__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11906__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07139_ _06755_ _06757_ _05658_ _06758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07586__A2 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10150_ _00358_ _02874_ _02955_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__13659__A2 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10081_ net63 _06691_ _02608_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07625__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13899__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07889__A3 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13840_ _00171_ clknet_leaf_51_clk DDS_Stage.xPoints_Generator1.RegP\[-8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_11_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13771_ _00106_ clknet_leaf_11_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10983_ _03822_ _03823_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12722_ _05599_ _05600_ _05601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10645__A2 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11842__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07360__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_26_clk_I clknet_3_7__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12653_ _05465_ _05525_ _05526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_155_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13595__A1 _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11604_ net54 _02051_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12584_ _05448_ _05449_ _05450_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09263__A2 _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07274__A1 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11535_ _04302_ _04376_ _04377_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07274__B2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11466_ _04277_ _04278_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07026__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13205_ _06121_ _06123_ _06124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10417_ _03227_ _03235_ _03294_ _03295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11397_ _04232_ _04238_ _04239_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_104_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08774__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13136_ _06047_ _06048_ _06049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10348_ _03138_ _03226_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__10581__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13067_ _05974_ _05975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_146_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10279_ _03052_ _03157_ _03158_ _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12018_ _04801_ net99 _04860_ _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11833__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07490_ _06703_ _00496_ _05182_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_66_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13586__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09160_ _02049_ _02050_ _02052_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_146_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ _01010_ _01011_ _01012_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_72_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13814__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09091_ _01896_ _01910_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11061__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08042_ _00938_ _00939_ _00941_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10644__B _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07812__I0 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09993_ _02872_ _02875_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_110_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08944_ _00398_ _06598_ _06618_ _00394_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09309__A3 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13510__B2 _06131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10324__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08875_ _01622_ _01684_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07826_ _05280_ _00398_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07757_ _00694_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10627__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-3\] _00652_ _00395_ _00653_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09427_ _02238_ _02316_ _00395_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09358_ _02179_ _02180_ _02247_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08309_ _01206_ _01210_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__13805__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07256__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09289_ _00376_ _06674_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11320_ _04076_ _04089_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07008__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11251_ _04076_ _04089_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10202_ _03080_ _03082_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_120_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11182_ _03956_ _04023_ _04024_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10133_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-7\] _03014_ _02935_ _03015_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08508__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13501__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10064_ _02867_ _02889_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_141_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10330__A4 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13823_ _00154_ clknet_leaf_68_clk DDS_Stage.xPoints_Generator1.RegF\[-10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13754_ _00089_ clknet_leaf_62_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11815__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11815__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10966_ _00393_ _02236_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09484__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12705_ _03189_ _00378_ _05582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13685_ _00020_ clknet_leaf_0_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10897_ _05387_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-22\] _03764_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07103__B _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12636_ _05394_ _05403_ _05506_ _05508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07247__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12567_ _05362_ _05432_ _05433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_124_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11518_ _00354_ _02499_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12498_ _05282_ _05348_ _05355_ _05358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_152_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11449_ _04259_ _04263_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10929__I0 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10554__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13119_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-8\] _05932_ _06032_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06990_ _06629_ _06630_ _06631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10306__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08660_ _06637_ _00376_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07611_ _00577_ DDS_Stage.xPoints_Generator1.CosNew\[-14\] _05182_ _00586_ _00587_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08591_ net73 _06659_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07542_ _05658_ _05529_ _00441_ _00443_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_72_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07473_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-12\] _00483_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07486__A1 _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09212_ _02028_ _02029_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_147_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09227__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07238__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09143_ net60 _06685_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12782__A2 _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09074_ _01959_ _01966_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08025_ _00878_ _00926_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07410__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09976_ _00370_ _06730_ _02829_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08927_ _01818_ _01821_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09163__A1 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08858_ _01751_ _01752_ _01753_ _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_93_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07809_ _00720_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08789_ _01685_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_123_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10820_ _03654_ _03658_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07477__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11273__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07477__B2 _06787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10751_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[1\] _03617_ _03623_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[2\]
+ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_36_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13470_ _06321_ _06327_ _06410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10682_ _05280_ _03556_ _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12421_ _05272_ _05273_ _05274_ _05275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11025__A2 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12352_ _05197_ _05198_ _05200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_22_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11303_ _04141_ _04145_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_132_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12283_ _04955_ _04956_ _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08729__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12525__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11234_ _04058_ _04059_ _04060_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07593__B _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07401__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11165_ _04005_ _04006_ _04007_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_140_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07952__A2 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10116_ _02995_ _02997_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11096_ _03906_ _03937_ _03938_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10047_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-9\] _02851_ _02848_ _02930_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_89_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_42_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold80 net168 net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold91 _05291_ net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_89_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13806_ _00137_ net36 clknet_leaf_73_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_86_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11998_ _04148_ _04156_ _04841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09457__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13737_ _00072_ net36 clknet_leaf_13_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_129_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11264__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10949_ _03790_ _03791_ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_70_clk clknet_3_0__leaf_clk clknet_leaf_70_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11803__A4 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13668_ _00003_ clknet_leaf_58_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-22\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08680__A3 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12213__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11016__A2 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12619_ _05399_ _05487_ _05488_ _05489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13599_ _06544_ _06547_ _06548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12516__A2 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08196__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09393__A1 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09830_ _02617_ _02714_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_74_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07943__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09761_ _02542_ _02645_ _02646_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06973_ _05919_ _06613_ _06615_ _06616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08712_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[4\] _01610_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09692_ _02578_ _02496_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer12 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-3\] net64 vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xrebuffer23 _00366_ net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08643_ _01458_ _01472_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xrebuffer34 net96 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
Xrebuffer45 _00362_ net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_77_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08574_ _01458_ _01472_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07459__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07525_ _05658_ _06651_ _06733_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09999__A3 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_61_clk clknet_3_1__leaf_clk clknet_leaf_61_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_147_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__A2 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07456_ _05409_ _06734_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07387_ DDS_Stage.xPoints_Generator1.CosNew\[-4\] DDS_Stage.xPoints_Generator1.RegP\[-4\]
+ _00402_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08959__A1 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09126_ _01924_ _02017_ _02018_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10766__A1 _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11963__B1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09057_ _01775_ _01949_ _01950_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_115_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08008_ _00394_ _05398_ _00844_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_60_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13180__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09959_ _02659_ _02663_ _02755_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09136__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12970_ _05763_ _05769_ _05868_ _05869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11921_ _04761_ _04763_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12691__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11494__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12691__B2 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11852_ _04666_ _04667_ _04653_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_129_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10803_ _03627_ _03675_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12443__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11783_ net66 _01693_ _01610_ net54 _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_68_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_52_clk clknet_3_1__leaf_clk clknet_leaf_52_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_45_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13522_ _06411_ _06429_ _06465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10734_ _03606_ _03607_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13453_ _06388_ _06390_ _06391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07870__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10665_ _03538_ _03539_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_12_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07870__B2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12404_ _05254_ _05255_ _05257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13384_ _06236_ _06255_ _06317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10596_ _03468_ _03471_ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_140_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12335_ _05151_ _05150_ _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_133_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07808__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12266_ _05055_ _05059_ _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13171__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11217_ _00365_ _02854_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12197_ _04366_ _05038_ _05039_ _05040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_50_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11148_ net84 _03485_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09127__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11079_ _03899_ _03920_ _03921_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09678__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11237__A2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08102__A2 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_43_clk clknet_3_4__leaf_clk clknet_leaf_43_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07310_ _06059_ _00358_ _00360_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08290_ _01179_ _01191_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_128_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10996__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07241_ _05409_ _06720_ _06774_ _06480_ _06146_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07172_ _06785_ _06786_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07718__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08169__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09905__A3 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09813_ net91 _06730_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11712__A3 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10920__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09744_ _00376_ _06701_ _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06956_ _05691_ _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__09669__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09675_ _02512_ _02561_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_38_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06887_ _05420_ _05474_ _05734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08626_ _05280_ _01524_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_120_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ _01395_ _01398_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_34_clk clknet_3_5__leaf_clk clknet_leaf_34_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07508_ _06146_ _05897_ _05182_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08488_ _01373_ _01387_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10987__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07439_ _05387_ _00449_ _00454_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12728__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10450_ _03324_ _03327_ _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_116_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09109_ _01998_ _02001_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11400__A2 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-5\] _03185_ _03183_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-4\]
+ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12120_ _04960_ _04962_ _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_107_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09357__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12051_ _00369_ _02409_ _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11164__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07907__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11002_ _03842_ _03844_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12953_ _05741_ _05821_ _05851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11904_ _04746_ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_116_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12884_ _05770_ _05775_ _05776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11835_ _04677_ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold90_I LoadP vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08096__A1 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11766_ _04601_ _04607_ _04608_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13505_ _06375_ _06377_ _06437_ _06446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10717_ _03585_ _03590_ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07843__A1 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07843__B2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11697_ _04539_ _04537_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_71_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12719__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13436_ _05387_ _06371_ _06372_ _06374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_10648_ _03453_ _03454_ _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_125_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer3 _02489_ net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13367_ _06289_ _06299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_125_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10579_ _03388_ _03453_ _03454_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_106_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07538__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12318_ _05140_ _05144_ _05161_ _05162_ _05163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__07071__A2 _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13298_ _06180_ _06181_ _06224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13144__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12249_ _05041_ _05044_ _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_149_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07790_ DDS_Stage.xPoints_Generator1.RegFrequency\[-4\] DDS_Stage.xPoints_Generator1.RegF\[-4\]
+ _00402_ _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_147_Right_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_134_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08859__B1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09460_ _02346_ _02347_ _02348_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_64_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08411_ _00869_ _00928_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_114_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09391_ _00357_ _06708_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_clk clknet_3_6__leaf_clk clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08087__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08342_ _01214_ _01230_ _01240_ _01243_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_46_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09823__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08273_ _01078_ _01174_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11630__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07224_ _05409_ _05485_ _05594_ _06830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_14_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09587__A1 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07155_ _05409_ _06732_ _06772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07086_ _06243_ _06711_ _06712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07062__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13135__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11146__A1 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08011__A1 _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12894__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08562__A2 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07988_ _00856_ _00861_ _00889_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09727_ _02526_ _02527_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06939_ _06265_ _06276_ _06287_ _06297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12646__A1 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09658_ _02438_ _02543_ _02544_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08609_ _01507_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09589_ _02469_ _02476_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11620_ _04460_ _04461_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10557__B net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09814__A2 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07825__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11551_ _00381_ _01693_ _01610_ _00384_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_107_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08093__A4 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _03305_ _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_133_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11482_ _04276_ _04281_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10975__A4 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13221_ _06136_ _06137_ _06140_ _06141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10433_ _03310_ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11385__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13152_ _05969_ _06064_ _06065_ _06066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_21_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08250__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10364_ _03139_ _03140_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12103_ _00381_ _01956_ _01794_ _00384_ _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13083_ _05915_ _05916_ _05992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10295_ _02141_ _02142_ _03174_ _02140_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_12034_ _04876_ _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_53_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11688__A2 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09750__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07093__S _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12637__A1 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12936_ _05830_ _05832_ _05834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12867_ _05663_ _05667_ _05758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_75_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11818_ net66 _01693_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13062__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12798_ _03340_ _00375_ _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11749_ _04589_ _04591_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13419_ _06333_ _06354_ _06355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13365__A2 _06295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08960_ _01852_ _01853_ _01854_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_110_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5_clk clknet_3_6__leaf_clk clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07911_ _06642_ _00352_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12876__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08891_ _01785_ _01786_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-21\] _01787_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11679__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07842_ _05864_ _05833_ _00388_ _00385_ _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_120_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07773_ _00702_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclone8 net76 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_16
X_09512_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-14\] _02400_ _02401_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10103__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09443_ _02260_ _02261_ _02331_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09374_ _02187_ _02188_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_136_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08325_ _01199_ _01211_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10406__A3 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08256_ net58 _00355_ _05833_ _05398_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_145_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07207_ _06232_ _05431_ _05658_ _06816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_115_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08187_ _01087_ _01088_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09024__A3 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11906__A3 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07138_ _06469_ _06756_ _06757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07035__A2 _06668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07069_ _06059_ _06695_ _06697_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11119__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10080_ net63 _06691_ _02608_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07889__A4 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13770_ _00105_ clknet_leaf_11_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_126_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10982_ _00369_ _02854_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12721_ _02854_ _00390_ _05600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10645__A3 _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11842__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12652_ _05502_ _05524_ _05525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_127_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11603_ _04443_ _04444_ _04445_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13595__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12583_ _05280_ net27 _05450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11534_ _04303_ _04304_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_92_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11465_ _04277_ _04278_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07596__B _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11358__A1 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold53_I FreqPhase[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13204_ _06122_ _06037_ _06123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10416_ _03230_ _03293_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08223__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07026__A2 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11396_ net66 net54 _02236_ _02153_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_150_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08774__A2 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09971__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13135_ _02940_ _00397_ _05989_ _06048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10347_ _03224_ _03225_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07816__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13066_ _05968_ _05972_ _05974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_146_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10278_ _03055_ _03069_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09723__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12017_ _04846_ _04858_ _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12919_ _05809_ _05814_ _05815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_66_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11833__A2 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13899_ _00230_ net36 clknet_leaf_18_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[21\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_66_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10892__I0 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-24\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13586__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08110_ net73 _06308_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08462__A1 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09090_ _01896_ _01910_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11061__A3 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08041_ _06598_ _00370_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10021__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09992_ _02779_ _02873_ _02874_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_86_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07726__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08943_ _01751_ _01836_ _01837_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_86_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09309__A4 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08874_ _01704_ _01706_ _01769_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07825_ _06059_ _00573_ _00728_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13750__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ net106 DDS_Stage.xPoints_Generator1.RegP\[-6\] _00684_ _00694_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07687_ DDS_Stage.xPoints_Generator1.CosNew\[-3\] _00651_ _00577_ _00652_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09426_ _02313_ _02315_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_48_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09357_ _00373_ _06679_ _02181_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_34_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ _01208_ _01209_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09288_ _00379_ _06672_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10835__B _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10260__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08239_ _01097_ _01117_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07008__A2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11250_ _04091_ _04092_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12001__A2 _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09402__B1 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10201_ _03081_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11181_ _03957_ _03958_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10132_ _02926_ _02928_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_128_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08508__A2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13501__A2 _06441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10063_ _02913_ _02921_ _02944_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13741__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07192__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13822_ _00153_ clknet_leaf_69_clk DDS_Stage.xPoints_Generator1.RegF\[-11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07319__I0 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13265__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07371__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13753_ _00088_ clknet_leaf_59_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11815__A2 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10965_ _00390_ _02238_ _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12704_ _05479_ _05481_ _05580_ _05581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13684_ _00019_ clknet_leaf_0_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10896_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-22\] _03763_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_38_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11028__B1 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12635_ _05397_ _05402_ _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11579__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_139_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12566_ _05430_ _05369_ _05432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_156_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11517_ _04299_ _04358_ _04359_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12497_ _05356_ _05282_ _05339_ _05344_ _05357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_103_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11448_ _04270_ _04283_ _04290_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11379_ _04208_ _04220_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10554__A2 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13118_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-8\] _05932_ _06031_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13049_ _00369_ _03679_ _05955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13732__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07610_ _00577_ _00585_ _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08590_ _01410_ _01487_ _01488_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13256__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_72_clk_I clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06930__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07541_ _05778_ _06721_ _06373_ _05658_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_89_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07472_ _06799_ _00308_ _00481_ _05658_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09211_ _02028_ _02029_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_91_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10490__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09142_ net61 _06679_ _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13799__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10242__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ _01963_ _01964_ _01965_ _01783_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_142_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_10_clk_I clknet_3_3__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08024_ _00907_ _00925_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_79_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09975_ _02826_ _02828_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08926_ _01819_ _01820_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09163__A2 _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08857_ net96 _06618_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07174__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13723__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07808_ _00370_ DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[21\] _00395_ _00720_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08788_ _01619_ _01622_ _01684_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06921__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07739_ _00685_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10750_ _03609_ _03615_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07204__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07477__A2 _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ _02200_ _02298_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10681_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[27\] _03556_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_47_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12420_ _05257_ _05271_ _05260_ _05274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_35_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07229__A2 _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12351_ _05198_ _05197_ _05199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_63_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06988__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11981__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11302_ _04144_ _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_133_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12282_ _04955_ _04956_ _05125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_120_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08729__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11233_ _04057_ _04065_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11164_ _03018_ _00372_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10115_ _02897_ _02898_ _02996_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11095_ net86 net83 _03416_ _03340_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10046_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-7\] _02926_ _02928_ _02929_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__07165__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold70 net164 net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold81 net167 net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold92 Enable net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__13238__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06912__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13805_ _00136_ net36 clknet_leaf_70_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11997_ _04819_ _04826_ _04839_ _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10948_ _00393_ _02238_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13736_ _00071_ net36 clknet_leaf_15_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__07712__I0 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10879_ _03747_ _03749_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_144_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13667_ _00002_ clknet_leaf_62_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-23\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_14_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08680__A4 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12618_ _05400_ _05401_ _05488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_143_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13598_ _06545_ _06546_ _06547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12213__A2 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10224__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12549_ net135 _00393_ _05413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06979__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09393__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13953__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09760_ _02545_ _02559_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06972_ _05713_ _06614_ _06615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08711_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-22\] _01529_ _01608_ _01609_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09691_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-13\] _02319_ _02393_ _02578_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__07156__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08642_ _01450_ _01538_ _01539_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xrebuffer13 _05149_ net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer24 _00362_ net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__06903__A1 _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer35 _04859_ net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xrebuffer46 _05445_ net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_1
XFILLER_0_95_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08573_ _01463_ _01471_ _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08105__B1 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07524_ _00419_ _00523_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10463__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07455_ _05387_ _00463_ _00464_ _00467_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_92_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07386_ _00413_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09125_ net137 net96 _06633_ _06696_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08959__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11963__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11963__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09056_ _01863_ _01866_ _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_114_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09908__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08007_ _00830_ _00835_ _00908_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_41_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11715__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13944__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09958_ _02841_ _02753_ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09136__A2 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08909_ _01721_ _01735_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_99_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09889_ _02693_ _02706_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11920_ _04760_ _04762_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12691__A2 _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11851_ _04676_ _04692_ _04693_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_79_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10802_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[3\] _03674_ _03675_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11782_ net70 _01524_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_103_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12443__A2 _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10733_ _03491_ _03536_ _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13521_ net147 _00397_ _06415_ _06464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_83_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13452_ _06337_ _06338_ _06389_ _06390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10664_ _03487_ _03489_ _03537_ _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_11_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07870__A2 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12403_ _05254_ _05255_ _05256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13383_ _06314_ _06315_ _06316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_152_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10595_ _03355_ _03469_ _03470_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12334_ _05152_ _04387_ _05179_ _04388_ _04408_ _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_50_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12265_ _05106_ _05107_ _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11216_ _00361_ _02938_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12196_ _04367_ _04368_ _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13935__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11147_ _03556_ _00351_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09127__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11078_ _03900_ _03901_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_10029_ _02890_ _02911_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_76_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11237__A3 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13719_ _00054_ clknet_leaf_13_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07310__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10996__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07240_ _05658_ _06698_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12198__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07171_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-20\] _06786_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09063__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11945__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13926__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ net73 _06742_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11712__A4 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07734__S _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06955_ _05409_ _06458_ _06469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09743_ _00379_ _06696_ _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07129__A1 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09674_ _02540_ _02560_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_38_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06886_ _05691_ _05713_ _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_27_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[3\] _01524_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_87_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08556_ _01378_ _01386_ _01454_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09826__B1 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07507_ _06726_ _06806_ _05658_ _05474_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_147_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08487_ _01378_ _01386_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10987__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07438_ _05387_ _00453_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07369_ DDS_Stage.xPoints_Generator1.CosNew\[-13\] DDS_Stage.xPoints_Generator1.RegP\[-13\]
+ _00402_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09108_ _01999_ _02000_ _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_131_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10380_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-4\] _03183_ _03259_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09039_ net60 _06679_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_131_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12050_ _04888_ _04892_ _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09357__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13917__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11001_ _03843_ _03793_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__11164__A2 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12113__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12952_ _05743_ _05849_ _05850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11903_ _04743_ _04744_ _04745_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10675__B2 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12883_ _05774_ _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11834_ _00361_ _01249_ _01247_ _00365_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_56_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07599__B _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11765_ _04603_ _04604_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08096__A2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10716_ _03388_ _03519_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold83_I rst vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13504_ _06365_ _06444_ _06438_ _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__07843__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11696_ _00381_ _01247_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10647_ _03453_ _03454_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13435_ _06365_ _06370_ _06372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_141_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer4 _01328_ net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_23_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13366_ _05822_ net22 _06298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10578_ _00385_ _06744_ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12317_ _05158_ _05159_ _05162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13297_ _06222_ _06223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_107_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12248_ _05089_ _05090_ _05091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13908__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12179_ _00381_ _00384_ _01794_ _01792_ _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__12104__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08859__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08859__B2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07531__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08410_ _00869_ _00928_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09390_ _02208_ _02278_ _02279_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08341_ _01241_ _01242_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_47_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08087__A2 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08272_ _01078_ _01079_ _01081_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11091__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11630__A3 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07223_ _05387_ _06824_ _06829_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11918__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07154_ _05822_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-22\] _06771_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09587__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07085_ _05420_ _05669_ _05409_ _06711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_2_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_113_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11146__A2 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08011__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12894__A2 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07987_ _00851_ _00855_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_89_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09726_ _02597_ _02611_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06938_ _05658_ _06265_ _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12646__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06869_ _05518_ _05529_ _05540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09657_ _02441_ _02444_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08608_ _01437_ _01506_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09588_ _02474_ _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10409__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08539_ _01358_ _01359_ _01357_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09275__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11550_ _04310_ _04318_ _04392_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11082__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10501_ _03362_ _03377_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11481_ _04211_ _04219_ _04323_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_18_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13220_ _06083_ _06138_ _06139_ _06140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_107_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10432_ _03138_ _03309_ _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07639__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12031__B1 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11385__A2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13151_ _05970_ _05971_ _06065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10363_ _03134_ _03240_ _03241_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08250__A2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12102_ _00387_ _01792_ _04945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13082_ _05915_ _05916_ _05991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10294_ _02225_ _02226_ _02490_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_103_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12033_ _04873_ _04874_ _04875_ _04876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_53_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09750__A2 _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12637__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12935_ _05626_ _05831_ _05832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07513__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12866_ _05754_ _05755_ _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11817_ _04657_ _04658_ _04659_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12797_ _03266_ _00378_ _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13062__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11748_ _04416_ _04590_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11679_ _00369_ _01430_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13418_ _06335_ _06353_ _06354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_141_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13349_ _06269_ _06279_ _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07910_ _06637_ _00355_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08890_ _01613_ _01606_ _01687_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__12876__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07841_ _06179_ _00382_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07772_ DDS_Stage.xPoints_Generator1.RegFrequency\[-13\] DDS_Stage.xPoints_Generator1.RegF\[-13\]
+ _00402_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09511_ _02310_ _02312_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclone9 net75 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XANTENNA__07504__A1 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _00373_ _06685_ _02262_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_84_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09373_ _02259_ _02262_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08324_ _01199_ _01211_ _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11064__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12873__B _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ _00993_ _01156_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07206_ _05387_ _06811_ _06812_ _06815_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_15_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08186_ _00953_ _00961_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_115_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09024__A4 _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07137_ _05572_ _05485_ _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11906__A4 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07068_ _05822_ _06696_ _06697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11119__A2 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10878__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07207__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09709_ _02530_ _02538_ _02594_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_126_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10981_ _03822_ _03823_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_12720_ _02762_ _00393_ _05599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12651_ _05505_ _05508_ _05523_ _05524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_11602_ net66 net54 _02051_ _01956_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_65_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12582_ _05360_ _05447_ _05182_ _05449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11533_ _04303_ _04304_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_52_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07369__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11464_ _04293_ _04306_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_52_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11358__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10415_ _03234_ _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13203_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-7\] _06027_ _06122_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_104_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08223__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11395_ net66 _02236_ _02153_ net54 _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07026__A3 _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10346_ _03222_ _03223_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_13134_ _05987_ _05988_ _06047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09971__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07982__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13065_ _05969_ _05970_ _05971_ _05972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_40_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10277_ _03055_ _03069_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12016_ _04858_ _04846_ _04859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09723__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12918_ _05810_ _05812_ _05813_ _05814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_88_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11833__A3 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13898_ _00229_ net36 clknet_leaf_18_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[20\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_66_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10892__I1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-24\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12849_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-10\] _05736_ _05738_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11046__A1 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08462__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11061__A4 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08040_ _00940_ _00941_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10021__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09991_ net60 _06744_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07973__A1 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08942_ _01752_ _01753_ _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_110_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08873_ _01714_ _01768_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_07824_ _05280_ _00394_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07742__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07755_ _00693_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_149_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11285__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07686_ DDS_Stage.xPoints_Generator1.RegFrequency\[-3\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-3\]
+ _00650_ _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09425_ _02314_ _02233_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13026__A2 _05840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09356_ _02174_ _02244_ _02245_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08307_ _00948_ _00969_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ _00373_ _06679_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ _01123_ _01136_ _01139_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10260__A2 _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12537__A1 _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08169_ _05864_ _00373_ _01042_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__07008__A3 _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09402__A1 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09402__B2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10200_ _00370_ _06744_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_152_Left_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11180_ _03957_ _03958_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10131_ _00506_ _03007_ _03012_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_24_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_128_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08508__A3 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ _02864_ _02912_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_128_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07652__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13821_ _00152_ clknet_leaf_72_clk DDS_Stage.xPoints_Generator1.RegF\[-12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_141_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09469__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07319__I1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13265__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13752_ _00087_ net36 clknet_leaf_43_clk DDS_Stage.xPoints_Generator1.CosNew\[-1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_134_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10964_ _00397_ _02153_ _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12703_ _05480_ _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_48_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13683_ _00018_ clknet_leaf_3_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10895_ _05822_ _06765_ _03762_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_48_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11028__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11028__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12634_ _05416_ _05425_ _05504_ _05505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11579__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12565_ _05372_ _05429_ _05430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_156_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11516_ net86 net83 _02499_ _02409_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_110_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12496_ _03773_ _05279_ _05356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_80_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11447_ _04256_ _04269_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_123_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11378_ _04208_ _04220_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07955__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10329_ _00398_ _06701_ _06708_ _00394_ _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13117_ _06029_ _06030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13048_ _05873_ _05879_ _05953_ _05954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13256__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07540_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[1\] _00537_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _05409_ _05442_ _05875_ _00480_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_88_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09210_ _02020_ _02021_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_17_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09141_ net73 _06691_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12767__A1 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10242__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09072_ _01787_ _01781_ _01868_ _01952_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_86_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12519__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08023_ _00909_ _00924_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_79_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09974_ _02766_ _02833_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08925_ _06654_ _00376_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08856_ net138 _06685_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07807_ _00719_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08787_ _01630_ _01683_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_54_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06921__A2 _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07738_ net2 DDS_Stage.xPoints_Generator1.RegP\[-15\] _00684_ _00685_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07669_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-6\] DDS_Stage.xPoints_Generator1.RegFrequency\[-6\]
+ _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09408_ _02294_ _02297_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10680_ _05182_ _03554_ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12758__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09339_ _00459_ _02144_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07220__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12350_ _05180_ _05181_ _05178_ _05198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_62_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06988__A2 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11981__A2 _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11301_ _04046_ _04142_ _04143_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_12281_ _05110_ _05114_ _05123_ _05124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_15_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11232_ _04051_ _04069_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11163_ _00375_ _02940_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10114_ _00373_ _06730_ _02899_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_11094_ net86 _03416_ _03340_ net83 _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10045_ _02838_ _02846_ _02927_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xhold60 net12 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__08362__A1 _06523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold71 net163 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold82 net171 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_89_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13238__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06912__A2 _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13804_ _00135_ net36 clknet_leaf_63_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_11996_ _04822_ _04825_ _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13735_ _00070_ net36 clknet_leaf_16_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_63_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10947_ _00390_ _02409_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13666_ _00001_ clknet_leaf_61_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-24\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10878_ _03311_ _03653_ _03748_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_155_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12617_ _05400_ _05401_ _05487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08417__A2 _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13597_ _00381_ _00384_ _03727_ _06546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_115_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12548_ _02499_ _00397_ _05412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06979__A2 _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12479_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-16\] _05338_ _05339_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_123_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06971_ _05550_ _05778_ _06614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08710_ _01606_ _01607_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11488__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09690_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-13\] _02394_ _02495_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-12\]
+ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_08641_ _01452_ _01503_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10160__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer14 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-14\] net88 vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06903__A2 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer25 _05740_ net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer47 _00366_ net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer58 _00778_ net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_08572_ _01466_ _01470_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08105__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12988__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08105__B2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07523_ _05940_ _06622_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07454_ _05182_ _00466_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10463__A2 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07385_ DDS_Stage.xPoints_Generator1.CosNew\[-5\] DDS_Stage.xPoints_Generator1.RegP\[-5\]
+ _00402_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clone13_I net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11412__A1 _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09124_ net96 _06633_ _06696_ net137 _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_60_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11963__A2 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09055_ _01797_ _01948_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07092__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08006_ _00827_ _00836_ _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09908__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11715__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08592__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09957_ _02749_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08908_ _01714_ _01768_ _01802_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09888_ _02691_ _02770_ _02771_ _02716_ _02736_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_08839_ _01726_ _01734_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11850_ _04690_ _04691_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07215__B _06822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10801_ _03667_ _03670_ _03673_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_0_131_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11781_ _04620_ _04622_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_103_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_103_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13520_ _06413_ _06414_ _06463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_45_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10732_ _03494_ _03535_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13451_ _03340_ _00397_ _06339_ _06389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13880__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10663_ _03487_ _03489_ _03537_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_11_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12402_ _04168_ _04146_ _05255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_136_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11403__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10594_ _03358_ _03404_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13382_ _06309_ _06310_ _06313_ _06315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_152_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07083__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12333_ _04371_ _04385_ _05179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13156__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07377__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_71_clk_I clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12264_ _04988_ _05001_ _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11215_ _00369_ _02762_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12195_ _04367_ _04368_ _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11146_ _00359_ _03416_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10390__A1 _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11077_ _03900_ _03901_ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07138__A2 _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ _02892_ _02895_ _02910_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_37_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_19_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06897__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11979_ _04811_ _04820_ _04821_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11237__A4 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11642__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13718_ _00053_ clknet_leaf_21_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07310__A2 _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_24_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13871__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13649_ _06594_ _06601_ _06602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_144_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13395__A1 _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12198__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ _06783_ _06784_ _05182_ _06785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_82_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09063__A2 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11945__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07074__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_39_clk_I clknet_3_5__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09811_ _02601_ _02694_ _02695_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10381__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09742_ _00373_ _06708_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06954_ _05572_ _05463_ _06458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09673_ _02542_ _02545_ _02559_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06885_ _05409_ _05702_ _05713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_38_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08624_ _01435_ _01521_ _05182_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06888__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07750__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08555_ _01381_ _01453_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09826__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09826__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13622__A2 _06563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07506_ _05387_ _00506_ _00509_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08486_ _01381_ _01385_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_65_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13862__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07437_ _06698_ _00450_ _00452_ _05658_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13386__A1 _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07368_ _00404_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07065__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09107_ _06664_ _00376_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07299_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-15\] _00352_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_115_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09038_ net92 _06674_ _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10747__I0 _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11000_ _00397_ _02236_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12113__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12951_ _05820_ _05849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11902_ _00381_ _00384_ _02153_ _02051_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_12882_ _05771_ _05772_ _05773_ _05774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07660__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11833_ _00361_ _00365_ _01249_ _01247_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__09817__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11624__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11764_ _04603_ _04604_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13503_ _06210_ _06294_ _06444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10715_ _03437_ _03587_ _03588_ _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13853__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11695_ _00381_ _01247_ _04537_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_138_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13377__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold76_I LoadF vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13434_ _06365_ _06370_ _06371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10646_ _03519_ _03520_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_153_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07056__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer5 _05199_ net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_13365_ _05822_ _06295_ _06296_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10577_ _00388_ _06742_ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12316_ _05158_ _05159_ _05161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13296_ _06219_ _06196_ _06220_ _06222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12247_ _04989_ _04997_ _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_39_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_71_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12178_ _00387_ _01693_ _05021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11129_ _03962_ _03963_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12104__A2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08859__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11863__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08340_ _01215_ _01225_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08087__A3 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08271_ _01074_ _01093_ _01172_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_74_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11091__A2 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11630__A4 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07222_ _05182_ _06825_ _06828_ _06829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_117_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ _05387_ _06765_ _06767_ _06770_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__11918__A2 _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12040__A1 _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07598__A2 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07084_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[0\] _06710_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08547__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13540__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10354__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__B1 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07986_ _00882_ _00887_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09725_ _02610_ _02605_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06937_ _06146_ _05529_ _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09656_ _02441_ _02444_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_2_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06868_ _05420_ _05474_ _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__10901__I0 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-20\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08607_ _01440_ _01505_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_78_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09587_ _00370_ _06701_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10409__A2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08538_ _01351_ _01421_ _01436_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09275__A2 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07286__A1 _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11082__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08469_ _01367_ _01271_ _01368_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10500_ _03368_ _03376_ _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11480_ _04214_ _04322_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10431_ _03307_ _03308_ _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12031__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12031__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07589__A2 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13150_ _05970_ _05971_ _06064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11385__A3 _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10362_ _03137_ _03151_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_33_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12101_ _04912_ _04940_ _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_103_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13081_ _05986_ _05989_ _05990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10293_ _03009_ _03172_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_130_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12032_ _00381_ _00384_ _02051_ _01956_ _04875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_109_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12934_ _05623_ _05723_ _05831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_137_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12865_ _05675_ _05689_ _05755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11816_ net66 net54 _01610_ _01524_ _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_12796_ _05570_ _05678_ _05679_ _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07277__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11747_ _04414_ _04415_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11678_ _00361_ _00365_ _01610_ _01524_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_40_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13417_ _06342_ _06352_ _06353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10629_ _03502_ _03503_ _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08226__B1 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08777__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13348_ _06273_ _06278_ _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_122_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13279_ _06200_ _06203_ _06204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07565__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08529__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07840_ _00738_ _00741_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10887__A2 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07771_ _00701_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09510_ _02150_ _02230_ _02231_ _02397_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XPHY_EDGE_ROW_56_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09441_ _02255_ _02328_ _02329_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_84_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09372_ _02260_ _02261_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _01219_ _01223_ _01224_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__13817__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07268__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11064__A2 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08254_ _01148_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07205_ _05182_ _06814_ _06815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_115_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08185_ _01054_ _01061_ _01086_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_65_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_99_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07136_ _06753_ _06754_ _06755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07067_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-3\] _06696_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07440__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10327__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09193__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07969_ _00824_ _00825_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_74_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09708_ _02516_ _02529_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10980_ _00365_ _02938_ _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09639_ net96 _06672_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07223__B _06829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12650_ _05513_ _05522_ _05523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_78_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13808__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11601_ net66 _02051_ _01956_ net54 _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12581_ _05360_ _05447_ _05448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07259__B2 _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11532_ _04372_ _04373_ _04374_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11463_ _04301_ _04305_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13202_ _06119_ _06120_ _06121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_10414_ _03276_ _03291_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07806__I0 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11394_ _04234_ _04235_ _04236_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08223__A3 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13133_ _05981_ _06044_ _06045_ _06046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07431__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10345_ _03222_ _03223_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07385__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07982__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13064_ _00372_ _03558_ _05971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10276_ _00373_ _06742_ _03059_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11515__B1 _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12015_ _04853_ _04857_ _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08931__A1 _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11818__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12917_ _03266_ _00381_ _05813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07498__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13897_ _00228_ net36 clknet_leaf_15_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[19\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_TAPCELL_ROW_66_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11833__A4 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12848_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-10\] _05736_ _05737_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11046__A2 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12779_ _05569_ _05574_ _05661_ _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10557__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09990_ net61 _06742_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07973__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08941_ _01752_ _01753_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_94_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08872_ _01716_ _01767_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_19_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07823_ _06059_ _00571_ _00727_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11809__A1 _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07754_ net108 DDS_Stage.xPoints_Generator1.RegP\[-7\] _00684_ _00693_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07489__A1 _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11285__A2 _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07685_ _00648_ _00649_ _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone43_I net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09424_ _00463_ _02228_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09355_ _02177_ _02191_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_63_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10245__B1 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08306_ _01185_ _01189_ _01207_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09286_ _02102_ _02175_ _02176_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_117_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08237_ _01137_ _01138_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12537__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08168_ _01040_ _01041_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_63_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09402__A2 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07119_ _05658_ _06740_ _06741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08099_ _00996_ _01000_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_24_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10130_ _02846_ _03009_ _03011_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10061_ _02919_ _02920_ _02942_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_128_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08508__A4 _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13820_ _00151_ clknet_leaf_71_clk DDS_Stage.xPoints_Generator1.RegF\[-13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_141_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09469__A2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13751_ _00086_ net36 clknet_leaf_42_clk DDS_Stage.xPoints_Generator1.CosNew\[-2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10963_ _03800_ _03805_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12702_ _05577_ _05578_ _05579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13682_ _00017_ clknet_leaf_0_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10894_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-23\] _03762_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11028__A2 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12633_ _05419_ _05503_ _05504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11579__A3 _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12564_ _05428_ _05405_ _05429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_156_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11515_ net86 _02499_ _02409_ net83 _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_135_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07400__C _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12495_ _03773_ _05279_ _05354_ _05355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_81_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11446_ _04285_ _04286_ _04288_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07404__A1 _06668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11377_ _04211_ _04219_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07955__A2 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13116_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-7\] _06027_ _06029_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10328_ _02704_ _03205_ _03206_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13047_ net70 _05765_ _05953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07128__B _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10259_ _00379_ _06738_ _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10711__A1 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13949_ _00280_ net101 clknet_leaf_26_clk net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_72_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_clk clknet_3_0__leaf_clk clknet_leaf_73_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07470_ _05409_ _00425_ _00479_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07891__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ _01931_ _02031_ _02032_ _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12767__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09071_ _00449_ _01961_ _01962_ _01953_ _01796_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_72_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12519__A2 _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08022_ _00910_ _00923_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_96_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09396__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09973_ _02769_ _02832_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08924_ _06649_ _00379_ _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08855_ _00355_ _06679_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10702__A1 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07806_ net61 DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[20\] _00395_ _00719_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08786_ _01632_ _01682_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_123_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12455__A1 _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07737_ _00683_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_123_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_64_clk clknet_3_1__leaf_clk clknet_leaf_64_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_149_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07668_ _00635_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09407_ _02295_ _02296_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_105_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07599_ _05387_ _00575_ _00576_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09338_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-15\] _02228_ _02229_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10769__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09269_ _02159_ _02072_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11300_ _04047_ _04048_ _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_132_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12280_ _05112_ _05113_ _05123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_133_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11231_ _04071_ _04073_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11162_ _04004_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09139__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10113_ _02892_ _02993_ _02994_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_140_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11093_ _03933_ _03934_ _03935_ _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_140_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10044_ _02834_ _02837_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12694__A1 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold50 net162 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_117_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold61 FreqPhase[2] net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08362__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold72 net169 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold83 rst net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_13803_ _00134_ net36 clknet_leaf_63_clk DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__12446__A1 _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11995_ _04832_ _04837_ _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_55_clk clknet_3_1__leaf_clk clknet_leaf_55_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13734_ _00069_ net36 clknet_leaf_23_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_EDGE_ROW_11_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10946_ _05822_ _00346_ _03789_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_63_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07873__A1 _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13665_ _00000_ clknet_leaf_61_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-25\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10877_ _03311_ _03585_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12616_ _05469_ _05484_ _05486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_14_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13596_ _00381_ _00384_ _03727_ _06545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07130__C _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12547_ _04000_ _04009_ _05410_ _05411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_41_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12478_ _05261_ _05337_ _05338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09378__A1 _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11429_ _04201_ _04202_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_20_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11185__A1 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10932__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06970_ _05409_ _05951_ _06613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07573__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11488__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08640_ _01452_ _01503_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10160__A2 _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer15 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-15\] net67 vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_83_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer26 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-13\] net78 vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12437__A1 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-20\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer37 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu1\[-3\] net136 vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_08571_ _01467_ _01468_ _01469_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__12437__B2 DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-21\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_clk clknet_3_4__leaf_clk clknet_leaf_46_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08105__A2 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-2\] _00522_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12988__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07453_ _05658_ _06656_ _00465_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_33_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07384_ _00412_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09123_ _01921_ _02014_ _02015_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07616__A1 DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07748__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09054_ _01863_ _01866_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_142_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08005_ _00880_ _00906_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09369__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09908__A3 _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11176__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08041__A1 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08592__A2 _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09956_ _02493_ _02839_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08907_ _01716_ _01767_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09887_ _02707_ _02715_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09541__A1 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08344__A2 _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08838_ _01729_ _01733_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08769_ _01587_ _01595_ _01665_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_leaf_37_clk clknet_3_6__leaf_clk clknet_leaf_37_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10800_ _03671_ _03672_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_11780_ _04620_ _04622_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_103_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10731_ _03560_ _03604_ _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_137_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07855__A1 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13450_ _06386_ _06387_ _06388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10662_ _03491_ _03536_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_125_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12401_ _04870_ _05252_ _05253_ _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_136_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07607__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11403__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13381_ _06309_ _06310_ _06313_ _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10593_ _03358_ _03404_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_36_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12332_ _05176_ _05177_ _05178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13156__A2 _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12263_ _05091_ _05099_ _05105_ _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11214_ _04052_ _04056_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08032__A1 _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12194_ _04382_ _05035_ _05036_ _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11145_ _03940_ _03986_ _03987_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_56_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07393__S _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12667__A1 _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11076_ _03890_ _03893_ _03891_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_10027_ _02900_ _02909_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07406__B _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06897__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_28_clk clknet_3_7__leaf_clk clknet_leaf_28_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11978_ net86 net83 _02938_ _02854_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_86_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__B _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10929_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-7\] DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-7\]
+ _05171_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13717_ _00052_ clknet_leaf_18_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11642__A2 _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07141__B _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13648_ _06597_ _06599_ _06600_ _06601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_30_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13579_ _06237_ _06476_ _06527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07074__A2 _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09810_ net61 net60 _06724_ _06730_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09741_ _02625_ _02626_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06953_ _05572_ _05680_ _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_20_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09672_ _02550_ _02558_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06884_ _05420_ _05463_ _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_38_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08623_ _01435_ _01521_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_38_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_19_clk clknet_3_7__leaf_clk clknet_leaf_19_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08554_ _01385_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09826__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07505_ _05182_ _00507_ _00508_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07837__A1 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11094__B1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08485_ _01382_ _01383_ _01384_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_65_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07436_ _05409_ _06092_ _00451_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07367_ DDS_Stage.xPoints_Generator1.CosNew\[-14\] DDS_Stage.xPoints_Generator1.RegP\[-14\]
+ _00402_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06890__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _06659_ _00379_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07065__A2 _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-15\] _00351_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_131_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09037_ _00357_ _06685_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09762__A1 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09939_ _02721_ _02735_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12950_ _05847_ _05845_ _05848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11901_ _00381_ _02153_ _02051_ _00384_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_99_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12881_ _00361_ _03679_ _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11832_ _04645_ _04674_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09817__A2 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07828__A1 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11763_ _04600_ _04605_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11624__A2 _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10714_ _03501_ _03504_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13502_ _06365_ _06438_ _06443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_83_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11694_ _04525_ _04530_ _04536_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13433_ _06131_ _06366_ _06369_ _06370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13377__A2 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10645_ _00388_ _00385_ _06744_ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_107_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11388__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold69_I FreqPhase[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13364_ _05280_ net21 _06296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10576_ _03388_ _03450_ _03451_ _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07300__I0 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12315_ _05069_ _05117_ _05159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13295_ _06145_ _06195_ _06220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_58_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12246_ _05078_ _05082_ _05088_ _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12177_ _04399_ _05018_ _05019_ _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11560__A1 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11128_ _03852_ _03969_ _03970_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12104__A3 _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11059_ _03899_ _03900_ _03901_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_64_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11863__A2 _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_86_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_103_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_153_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07819__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08087__A4 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08270_ net68 _01092_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07221_ _06826_ _06827_ _06828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07152_ _05182_ _06769_ _06770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12040__A2 _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07083_ _06059_ _06707_ _06709_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8_clk clknet_3_2__leaf_clk clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12879__A1 _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08547__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09744__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13540__A2 _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10354__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__B2 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07985_ _00885_ _00886_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09724_ _02606_ _02608_ _02609_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06936_ _05734_ _06221_ _06254_ _06265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09655_ _02456_ _02464_ _02541_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06867_ _05409_ _05507_ _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_2_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08606_ _01442_ _01504_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_96_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09586_ _02471_ _02473_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_70_clk_I clknet_3_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08537_ _01354_ _01420_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10409__A3 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08468_ _01262_ _01266_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08483__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11082__A3 _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07419_ _06624_ _00343_ _00437_ _05658_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_18_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08399_ _01274_ _01299_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_64_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10430_ _00379_ _00376_ _06744_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_21_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12031__A2 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11385__A4 _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ _03137_ _03151_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12100_ _04872_ _04942_ _04943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_14_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13080_ _05987_ _05988_ _05989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10292_ _03007_ _03091_ _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12031_ _00381_ _02051_ _01956_ _00384_ _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_148_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_23_clk_I clknet_3_6__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12933_ _05270_ _05439_ _05830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13047__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12864_ _05662_ _05674_ _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11815_ net66 _01610_ _01524_ net54 _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12795_ _05571_ _05573_ _05679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_139_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11746_ _04577_ _04581_ _04588_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08474__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11677_ _04519_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_43_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10628_ _00398_ _00394_ _06730_ _06738_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_13416_ _06346_ _06350_ _06352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08226__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08226__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13347_ _06274_ _06275_ _06277_ _06278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08777__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09974__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ _02704_ _03433_ _03434_ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13278_ _06201_ _06202_ _06203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12229_ net87 _02584_ _02499_ net84 _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_120_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07770_ DDS_Stage.xPoints_Generator1.RegFrequency\[-14\] DDS_Stage.xPoints_Generator1.RegF\[-14\]
+ _00402_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13286__A1 _06131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07581__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _02258_ _02272_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11049__B1 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09371_ _00376_ _06679_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08322_ _01221_ _01222_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07268__A2 _06125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08253_ _01146_ _01154_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07204_ _06646_ _06813_ _05658_ _06814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08184_ _01057_ _01060_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07135_ _06232_ _06458_ _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07756__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11772__A1 _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07066_ _05658_ _06694_ _06695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_113_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09717__A1 _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10327__A2 _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11524__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09193__A2 _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ _00837_ _00839_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10910__S _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06951__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06919_ _05420_ _06070_ _06081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09707_ _02540_ _02560_ _02592_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07899_ _00771_ _00799_ _00800_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08153__B1 _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09638_ _00355_ _06738_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07504__B _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09569_ _02380_ _02381_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11600_ net70 _01794_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12580_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-13\] _05446_ _05447_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_154_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11531_ _04314_ _04315_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11462_ _04302_ _04303_ _04304_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09405__B1 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13201_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-6\] _06118_ _06120_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10015__A1 _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10413_ _03282_ _03290_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11393_ _04229_ _04233_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08223__A4 _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13132_ _05985_ _06000_ _06045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_33_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07666__S _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10344_ _00376_ _06744_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13063_ _03556_ _00375_ _05970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10275_ _03057_ _03058_ _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__11515__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11515__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12014_ _04855_ _04856_ _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07195__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13744__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08931__A2 _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06942__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11818__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12916_ _03189_ _00384_ _05812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08695__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07498__A2 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09892__B1 _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13896_ _00227_ net36 clknet_leaf_18_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[18\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_57_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_66_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12847_ _05723_ _05726_ _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_61_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12778_ _05564_ _05660_ _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11451__B1 _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11729_ _04560_ _04565_ _04571_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10557__A2 _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ _01745_ _01746_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_94_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11506__A1 _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08871_ _01737_ _01766_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07186__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13735__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07822_ _05280_ net63 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07753_ _00692_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11809__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07684_ DDS_Stage.xPoints_Generator1.RegFrequency\[-4\] DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-4\]
+ _00644_ _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08686__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09423_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a1_in\[-14\] _02310_ _02312_ _02313_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__10493__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clone36_I DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[15\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09354_ _02177_ _02191_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10245__A1 _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08305_ _01187_ _01188_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10245__B2 _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09285_ _02105_ _02108_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07110__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08236_ _05833_ _00370_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09938__A1 _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08167_ _00986_ _01067_ _01068_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07118_ _06092_ _06622_ _06713_ _06740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08098_ _00997_ _00998_ _00999_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_3_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07049_ _06059_ _06678_ _06680_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _02941_ _02918_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13726__RN net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07177__A1 _06787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07218__C _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06924__A1 _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09469__A3 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13750_ _00085_ net36 clknet_leaf_45_clk DDS_Stage.xPoints_Generator1.CosNew\[-3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08677__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07234__B _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10962_ _03801_ _03804_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_12701_ _03018_ _00378_ _05497_ _05578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_97_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10893_ _03761_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13681_ _00016_ clknet_leaf_3_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a2_in\[-9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12632_ _05424_ _05503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12563_ _05408_ _05427_ _05428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__11579__A4 _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07101__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11514_ _04301_ _04305_ _04356_ _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_61_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12494_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[-15\] _05281_ _05354_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09929__A1 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11445_ _04253_ _04287_ _04284_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold51_I FreqPhase[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11376_ _04214_ _04218_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_156_Right_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10327_ net63 _06708_ net57 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_131_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13115_ _06015_ _06026_ _06027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07409__B _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13046_ _05949_ _05950_ _05952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09157__A2 _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ _00373_ _06744_ _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07168__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10189_ _03052_ _03055_ _03069_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__07144__B _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13948_ _00279_ net101 clknet_leaf_26_clk net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__08668__A1 _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13661__A1 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13879_ _00210_ net36 clknet_leaf_61_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.delay2.d_out\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__06983__B _06623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13413__A1 _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07891__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09093__A1 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11975__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09070_ _01961_ _01962_ _00449_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_71_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08021_ _00917_ _00922_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09396__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13956__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09972_ _05822_ _02853_ _02855_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08923_ _06659_ _00373_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07159__A1 _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12152__A1 _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08854_ _01670_ _01678_ _01749_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06906__A1 _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07805_ _00718_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08785_ _01653_ _01681_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07736_ net36 _05324_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08659__A1 _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07667_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-6\] _00634_ _00395_ _00635_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_105_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09406_ _06642_ _06649_ _00398_ _00394_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_105_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13404__A1 _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07598_ DDS_Stage.Block_Cosine.agu_1.agu_urgn_in\[-1\] _05182_ _00576_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_36_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09337_ _02156_ _02227_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_146_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11966__A1 _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09268_ _02070_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_138_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08219_ _01119_ _01120_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_44_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09199_ _06659_ _00382_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11718__A1 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11230_ _04037_ _04038_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07398__A1 _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13947__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11161_ _00378_ _02938_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09139__A2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ _02895_ _02910_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11092_ _00365_ _03189_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10043_ _02924_ _02925_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08898__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12694__A2 _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold51 FreqPhase[7] net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold62 net9 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold73 _05215_ net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold84 FreqPhase[13] net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_13802_ _00133_ net36 clknet_leaf_64_clk DDS_Stage.Block_Cosine.PolyRAM_1.delay1.d_in\[30\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__12446__A2 _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11994_ _04835_ _04836_ _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_86_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10457__A1 _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13733_ _00068_ net36 clknet_leaf_20_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.datax_argu2\[-5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_10945_ _05280_ DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.awire1\[1\] _03789_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13664_ _06146_ _05387_ _00576_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10876_ _03746_ _03710_ _03638_ _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07873__A2 _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12615_ _05478_ _05483_ _05484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13595_ _00387_ _03725_ _06544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12546_ _04003_ _04008_ _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12477_ _05336_ _05268_ _05273_ _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09378__A2 _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11428_ _04201_ _04202_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13938__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11185__A2 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11359_ _00372_ _01792_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07139__B _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10932__A2 _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13029_ _05848_ _05933_ _05934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10696__A1 _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07561__A1 _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10160__A3 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer16 _01076_ net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08570_ _00385_ _06598_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer27 _03342_ net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer49 _03416_ net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_88_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07521_ _05387_ _00517_ _00519_ _00521_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_88_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07452_ _05496_ _05713_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07383_ DDS_Stage.xPoints_Generator1.CosNew\[-6\] DDS_Stage.xPoints_Generator1.RegP\[-6\]
+ _00402_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09122_ _01923_ _01936_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09053_ _01943_ _01946_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_115_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08004_ _00888_ _00905_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__09369__A2 _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09908__A4 _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13929__RN net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11176__A2 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08041__A2 _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07764__S _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09955_ _02660_ _02574_ _02659_ _02755_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12125__A1 _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08906_ _01799_ _01800_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09886_ _02707_ _02715_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09541__A2 _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08837_ _01730_ _01731_ _01732_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__07552__A1 _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08768_ _01590_ _01594_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07719_ _00674_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08699_ _01581_ _01583_ _01596_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_68_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10730_ _03563_ _03603_ _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07855__A2 _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10661_ _03494_ _03535_ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12400_ _04863_ _04864_ _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_149_Left_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_11_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13380_ _06259_ _06311_ _06312_ _06313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_153_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10592_ _03419_ _03467_ _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__A1 _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12331_ _05170_ _05174_ _05177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12262_ _05089_ _05090_ _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11213_ _04053_ _04055_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12193_ _04379_ _04380_ _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08032__A2 _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 net30 Cos_Out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07674__S _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11144_ net86 net84 _03485_ _03416_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_56_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11075_ _03896_ _03916_ _03917_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10026_ _02907_ _02908_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07543__A1 _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09296__A1 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11977_ net86 _02938_ _02854_ net83 _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13716_ _00051_ clknet_leaf_17_clk DDS_Stage.Block_Cosine.PolyRAM_1.DataMac.a0_in\[-5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10928_ _03780_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13647_ _00397_ _03558_ _06600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10859_ _03592_ _03702_ _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13578_ _06478_ _06500_ _06525_ _06526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12529_ _05376_ _05390_ _05391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_140_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__A1 _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12107__A1 _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06952_ _06059_ _06405_ _06427_ _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09740_ _02443_ _02537_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

