`timescale 1ns / 1ps

module aguCosQI2_16b
#(	parameter DATA_WIDTH=16, 
	parameter ADDR_WIDTH=5, 
	parameter I_width =3, 
	parameter F_width=DATA_WIDTH-I_width
)
(	input agu_clock_in,
	input agu_reset_in,
	input agu_control_in,
	input signed [I_width-1 : -F_width] agu_urgn_in, 

	output [(ADDR_WIDTH-1):0] agu_address_coef_out,			
	output signed [I_width-1 : -F_width] agu_urgn_out
);
	
reg [(ADDR_WIDTH-1):0]		agu_address_coef_out;
reg [I_width-1 : -F_width]	agu_urgn_out;

always @(posedge agu_clock_in or negedge agu_reset_in) begin
	if (!agu_reset_in) begin
		agu_address_coef_out <= 0;
		agu_urgn_out <= 0;
	end

	else begin		
		if (agu_control_in) begin
			agu_urgn_out <= agu_urgn_in;

			casez (agu_urgn_in)
				16'b000001_?????????? : agu_address_coef_out <= 5'b0_0001;
				16'b000010_?????????? : agu_address_coef_out <= 5'b0_0010;
				16'b000011_?????????? : agu_address_coef_out <= 5'b0_0011;
				16'b000100_?????????? : agu_address_coef_out <= 5'b0_0100;
				16'b000101_?????????? : agu_address_coef_out <= 5'b0_0101;
				16'b000110_?????????? : agu_address_coef_out <= 5'b0_0110;
				16'b000111_?????????? : agu_address_coef_out <= 5'b0_0111;
				16'b001000_?????????? : agu_address_coef_out <= 5'b0_1000;
				16'b001001_?????????? : agu_address_coef_out <= 5'b0_1001;
				16'b001010_?????????? : agu_address_coef_out <= 5'b0_1010;
				16'b001011_?????????? : agu_address_coef_out <= 5'b0_1011;
				16'b001100_?????????? : agu_address_coef_out <= 5'b0_1100;
				16'b001101_?????????? : agu_address_coef_out <= 5'b0_1101;
				16'b001110_?????????? : agu_address_coef_out <= 5'b0_1110;
				16'b001111_?????????? : agu_address_coef_out <= 5'b0_1111;
				16'b010000_?????????? : agu_address_coef_out <= 5'b1_0000;
				16'b010001_?????????? : agu_address_coef_out <= 5'b1_0001;
				16'b010010_?????????? : agu_address_coef_out <= 5'b1_0010;
				16'b010011_?????????? : agu_address_coef_out <= 5'b1_0011;
				16'b010100_?????????? : agu_address_coef_out <= 5'b1_0100;
				16'b010101_?????????? : agu_address_coef_out <= 5'b1_0101;
				16'b010110_?????????? : agu_address_coef_out <= 5'b1_0110;
				16'b010111_?????????? : agu_address_coef_out <= 5'b1_0111;
				16'b011000_?????????? : agu_address_coef_out <= 5'b1_1000;
				16'b011001_?????????? : agu_address_coef_out <= 5'b1_1001;
				16'b011010_?????????? : agu_address_coef_out <= 5'b1_1010;
				16'b011011_?????????? : agu_address_coef_out <= 5'b1_1011;
				16'b011100_?????????? : agu_address_coef_out <= 5'b1_1100;
				16'b011101_?????????? : agu_address_coef_out <= 5'b1_1101;
				16'b011110_?????????? : agu_address_coef_out <= 5'b1_1110;
				16'b011111_?????????? : agu_address_coef_out <= 5'b1_1111;
				default : agu_address_coef_out <= 5'b0_0000;			 
			endcase														 
		end
	end	  
end 

endmodule  

